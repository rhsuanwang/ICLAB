`ifdef FUNC
`define LAT_MAX 20
`define LAT_MIN 1
`endif
`ifdef PERF
`define LAT_MAX 20
`define LAT_MIN 1
`endif

module pseudo_DRAM_data#(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=16, BURST_LEN=7) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface 
      // axi write address channel 
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [BURST_LEN-1:0]   awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------
   
      // axi write data channel 
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,
   
      // axi write response channel 
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master 
      input wire                  bready_s_inf,
      // -----------------------------
   
      // axi read address channel 
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [BURST_LEN-1:0]   arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------
   
      // axi read data channel 
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);
// Modify your "dat" in this directory path to initialized DRAM Value

parameter DRAM_p_r = "../00_TESTBED/DRAM/DRAM_data.dat";
// Modify DRAM_R_LAT           for Initial Read Data Latency, 
//        DRAM_W_LAT           for Initial Write Data Latency
//        MAX_WAIT_READY_CYCLE for control the Upperlimit time to wait Response Ready Signal
//
//        reg [7:0] DRMA_r [0:4*64*1024-1] is the storage element in this simulation model

parameter DRAM_R_LAT = 1, DRAM_W_LAT =1, MAX_WAIT_READY_CYCLE=300;
reg	[7:0]	DRAM_r	[0:8191];   // addr from 00000000 to 000203FF

integer dram_r_lat;
parameter LAT_MAX = `LAT_MAX;
parameter LAT_MIN = `LAT_MIN;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
CzUUnDspumJozn23NHO/AJQgR0Lj9Ze688saahOk+8kPJDHVjj8ovu+IHWByzgIc
oxM+lO4LC0yfECORZ25RMIiprG6vJAY2jXZ8++w8yvGzYHXgDV9mEAiIE8aw2Kfu
yx7nhk4iOHfoUhwB+1F1cI2sAB1h8WR8256qVcG/bFmktea+/7VDCg==
//pragma protect end_key_block
//pragma protect digest_block
+62RAhKwrrE40orUYRd+LVeUp6c=
//pragma protect end_digest_block
//pragma protect data_block
lyf3LyHHybO7XevA8ZmhnLCqAbenylS6JuZ16lZ4LaE2n1tg1/A3Lt2oyJ1mzbQt
34w+i+IQi/4z3Jojr+64XTo7G4BorPiZXS7gHW0rf1RL4CUKr0AES+CFpRTe9Jy3
78oM53wnWWboSq+l0ucqQltodSonemxXBW5lfAk3GU2MtV4OYChSo1/yrrAW/DFn
edxaeBfzcXTXNoXv/Pe8H5sFG3vSUr1FkAFZrf1J0vTlxlNYeNiPqmJ103wktL6r
jXFiszNy4QLcXCf35FIXN8/ghmfsl4iHnhpeQGxmWeJDFssgNb7Y2fr5bhOwV7cn
5bvQmC9yiKEpSMJPUWevmBAlDvYNUUWz6YmqoIu8xvtCTo5ie7Y2EEd4qDS0E0E7
72NTnjuADFyVh/vGR1WeEw5DussIigvslw7j8pwg1Y5dKE66PFLUv80X/bZ1MCDd
3PBbTDNnqMU4fxYo9eMpt2C+zhgm+zfEW/7b7tbeinjmpkftGVHySoAuerMO0ty+
oPjTMv7TI2VEYq4OcxmgPoom1oiM5Kh4f0Gsze4jToF6+1v+Y9mXiLEFbyRZfA+G
buDieY2+dbVfjEWxTkVJPoSCPKTB3iT+GcgHMgYiM9euFYfGzDVXrtsKzC7At85z
iRdqA+Ex5X3yZNJNQfyNX2rlFpfMpAr1zIXkp2Lj82s8zp75OuNDFPmMOMELHM1h
Ied+sDUzDaMsrm2s1DuUImR67z/7xk/vCzlSYjEupuFlKdDJ6qcwWLWyWg2Jg9O9
b1vAm2wTLezNrqs++tSgNq7FE3o/6e5Ch4EZxIGgvyGVru1GsOcoY9acqgzwRLie
auC31mEamLdJwc9tIgOrnh1xbW9pxSuwE0so2u7MOZAI9LrmW/+Kwfi0tBycCU7F
GsyY62rVPDdVdQv47Xh5Qkd2X8oXWLuzBb2IZ+y3kxJ2k6DrRMVyIKdz79YzE+29
cbiC6oEyuecOOZaFGlAAL4ZzaCpoeTbVi7g06gklf71g9MaG58o73XkXHco6fj9Y
hm9QE2RSJ27Xv20G6sqqdqklElE5kNOTifhwwd1D7W6KAjg1pTH1G2YswtQPy7/V
8d34hswopMuDpRJj7oLxi9oQnTbgbHg9STlCp81TzBYlgTL7ShDwXp7ijihn53jI
s4OfrpShjrAbXsQzdQZVoi5D73inZ9m0c+kqW70hMIyI0qrx8EsgUYSyJRwvQQu6
um/nRWe9h2Ul2cxeSGm+LkfxrkDubbGh0hvBqYdBs4BsxCYRCrE1fgVUCsJYFqlZ
7Zx1NKublIcmHJlSzlRd4AW0FBYu6FYbcoRSC/+JwKRENgtftnScSPhaZDeNG85L
BEU32ruBp+6gMmu0htlo5mUn/KCNay6j67u1ddP8igsBh7DasVBqfILTrR27MeRF
Jf5VroQa1TIRY2QWorCDGy22z7ulUvaSrguEyUIF2RpL1tOXXlMHlZiRQkiGZB4A
TjEvm1xoVGxq4h37cHYmI+4RrV5SRP0eKrul2/aCdZ2NOjpkAny8JAPqUymip5pd
8NDY3vLGp/4MkB3wRf0zNJ3TKBFykI/LvOYzl7JLkZVkoL30eJmogF4vlbrWuRs0
V1+kXlZwFWXtPURr5mGO9f/B9jOu625F+fquK5sTTuyYJo3+BCHsxHfC6i2LRTYF
CPsnfriYJtwwHmrTU+CeFZ6tfWckK7NNx9hLfCrFe5EkUiMblGQXEqtV86OtKIcb
k5dTQFJXKLGrcqoonzVAXlkgHl6NPscT6qWJ6qLAhCO7LX2iKOtThA5qIaQgS+Ph
rDb1W3tDa6oi6KjzgNmJ7OiG3n2Iy/EcIvzirfsGwJCp0h/B8CHMAq35rVbAtA+V
ZKae0y9hK3e8sxwW6w1kGSGyfSUnoiy48SKG/8742UZ3RksO6a/P8WavgUVrEOc3
IZVbHLVaGIpl7M+HVb0v20p6jp767O2PRQzlCojdpl7cr6XnDeHVBuKmsMgLieqf
UTS0lY6mMPSpXjOWNlEOp/Jb82IadIK1C7xntvEtaiG4zUJH17v8SZcvNJhHn/T8
sKjQt2o6nTmzTCR1S9FBg085w4PaQ87wBVb7CzM+zbmN4zQeT+P3a+diikPl2A3/
ihpgvOyBDvU5xhvBCT3HjLyS0rVwCk+gOzh/ZZc7udtQmYOiXbYH4ILBfGY9ZFZ8
V+PAGhzqRWxXuIwApArrKJ83esGXV23zocOLKzcgLU1nlWmThYuWhvjBy3RH2nTO
3VCwJFzbvzYCMILHHpFH+uWNGUUqRs7tEl2tj9MdUuLH2wilxCwfeG3poueLStk2
14sBGG0MyII69/SdV8iGdGdsGrzoEuTI9z+W9l0+TDmRMX618bTWJHj8p1MRvc9f
Lkx2S2wW2W8oOqpRDWMd6zgJ3S5ktU9VgJ9D/NEC66JZQrz1nkeN/PUo2VOIOmzw
y4+/6dSnSZlIfjQumqCoK2dSTN2tavadnc7YCIEo1PB82OdCydRQbHcDrRrlEUBr
XwcI8XCi5fNGig6DOmHO893v1dUsOhHAf249yOfcitvfNNfFUMCZJvECTDO1g/Rn
DB5CR7V18C67NU0+7m7c7yvcCiTJhvC5P5y6DhH2QGDfJalCt0XSbuVXtzZeuonB
IEQ86BOehDB+YiG4O0i5ZlqOVVkS9WejdxFockxj1OeWxJdCGaz5kKuuBljDSHvr
ViXyfaDMzqOnpYAAjpKvSSHAx044QIDJ1mLtkHr6B1pQNxU2tptJGIhVb2vahedu
ysWSN24d8ctKr7VC9hxS6uXYHLvhT2ZoWOg1KbJ0cXH0atS/uPdBz5KNgRlwLVYq
T+8b174XHPW3yWWynwE804y6EWtdH56wEbqbmZSdCCPTQnwvWP8OkOt3Y03GA06/
8vBLj5LaDqkgXNXDkfI6DzAAsRE/pQB0eZam1FMHRnt1CexuAlDE2AoRVgZFIIbk
MgPkL5dNfA39ZUime4QtKsCeHKO5J8gkI3/ujUMEX+dG3Gs4lunrakJUv+0rTjf+
Hl6AGNDVAbFLvYvdCi4ARrIQS9FjdpDVUH5Eu+wD792GzV2B+a6cSXWysvKz9YDG
L8QxZDB2+4UHKKfrVhMQ8P/RQqXOCoN62YketBZBCySa5t0Bb9n61MIdVHKwGaoI
Osuj0WyUpKKrBuZsjaUS6gPgJkbX3REzYv2iRhzs9y6H22NIwAUzkX3ZWQGLqD4w
fTtb6mOWDuyr1CtqVIEXLCKLn0XoLCK/YxkVWKf2bzFvglLR4kQfQdiQ1O/II7MD
dMR7NrKLYa22VGQybKqOoV7yBBrxFb6SSXZjwQy96ZGxzKBDfNFBgIMsH56o5Jo/
ymm4Ljk9YutgWnooAlYL1VoZQjh1PaMj6BtJErdLWxvKoc+6JkLQS1c990lRiLo3
I3/Gqq0rWydcR9tl3K93LZUyBzStmQDkJHwkzG1EulKDzoRUd2qN9c0tW8+hfsTa
tcq2Db4Sy5N4foZDQv2ZMb5ZXxACCq331uYm6Oe8r1CBSJYHIHEaGEUkBm8gaNUD
CwO8X00FAPiNEHoSq20HteXMuMXo01p2CmKOQhpYhOJGLnj1FqJkmyVsQ/qHAt9K
G5DhgbY3vcWRniRxoVA8oSgiAKR01N5KZvoCcec4/dGWzLl3OkETrBU0/gBK/k1J
djOu0towBNobP70MjxypS7uHTAtq2qiVhX0BrcYXkMosPiE/PRXwYn0vBSixet7q
dP6w7RykQc/OuDTSNdp4ThpX9aafThqzGA4kLgnGn3jC+Uo4wSi44CBfzbKGa1A1
h88ogAojOmely0J7hux6OiH07NG6NBpk0Zdx2DbVaA+TGRtVjLNA7/xNDBqMrtG4
7pW5zHBiey5mgT4ReKcmM/ss6Ny//2xLBScLSd1iAbyDZmRUoKyV/oHHWZIi0zZS
LjGZtIa6NXTCbwyN1HkU0sJGib/hdCaBKQIP/5JEd7X21kIsB+yNsj199GSB3bfT
pRuQ8FZeAouo9sAJruNM4BhC447x9ASG4axOXZuzEFo3rwEcmjioDmPyy2T3hf60
fHPRp2s0GfdVClsnJecBZtJKPZKMPOLW+FSlRhF5VJDmjYKS9DHePCSvLYFh1IWD
E6LxLYRMyg0F9eN480ER749vg3rzhaetD04YgUm9O4aBGXycK8JL+kgPntUDutk1
XBtjSMrrS6Tes1fDF4DN3FqUm5vz1yjjLquvSJhhCSW9Eh/Kan4XQsX53iSAcjok
yTeLJBZsGoZ109VXTMDT0vEH/nbsJx/XTBO/9RQuLJ2vZBFBjcGQLNVY24sA7KRU
bb+Lx8bt5aMgw51rusUT7yxzF35N1iweYF7rEZAlMKdtEodifcr3Ea/xvDCZG7ZY
9XGtfuu1uXcSEgk9yrknAYepJrGeVJenV0/BBnApmgg/gH4LE2ORbgw1GRTqDTgw
EM6g6DTIPd5osWcR4OzkEFJ2q6r9hQxdh5qkC9+Aun9ysCU2O+ARgxtq8MOBKudr
SASQLV/x3lrWkZBlpbkBcNA/rL0ezcs70y1gMM5lop++LSWu1sIfHTS8CZ0U4hDO
tjMY5rf6RSuMwqfu/ULHE3n7FdBnsJca8znGsZLu+V0DYNcoLkGzt45qGmRmrygq
Bh9dJof9ISyamIloU7G2VaBN115pgX4mwhdQtoH/uLR/7bcOaUqtckYS55giXDl6
vxHYJAN/BPIwMZLd3HvUgPqsJvZKFz/rGUUxJcJpRriRCv68MoBF0h/E+y3N9PTG
L/p2IU8EvnRy+R39UzQcgLikIe5AET5AmIlKlRUKyk5FKycUrR1gzLgXTXiTvxEX
6MOI7L+2ep3hjyQIrT7LKNHf9hAH3ZrNX7dUUrNeLEBQ42Ny55ud0pIoFxvzGIcu
zU84dlnuHi4nUA97gGbi9faMPNYmQAkxQ7kvvWyRVXljGaAFFd41pwvOGSsF58F/
AP8rq022ebNJ1d/BDP4pgjHq9xWGcvKMBne5DIlrN62IYMMiMtxz+Op2siH5DRGd
SO+5sqtqWMPW+Xo1cXhFdahJGybJ9NQJASziP1rYx5GjuGvcRCDRDxwaf9XHmW8l
ejIANsCWdkbdOmMYisTXN/D4Z3W0k73cT78Kq/MUEEGRi3pgg9C/SedMS99jbXv8
QB72C8a7Lhonm6jFT4ZGiI1MQopHNnKNDq4cD4nYQtUTFOW15FezRISsfa7vmLhb
zmMJQJ1NbuA6OyBgEHMzf1CaCQkyajaLU9YlmUIKmXS8fheujYmc6IHQf+cFOEDH
RIQU1kprTStEo4NWcWOwhdL6UbzOU2NTwxQEbFQWFp1GDG/72woiDfNh5G3UlkAM
v8HdnX52UBsiPwdgt5VNkrgWUk/qdeoSQ9pdO3QgigpPpptR3ellVUucrOphmeuj
vL90dq2S4yaCs7Apwn8c0nCfrlKWG2S0WhtCkiaafHcbWA2FFOl6GBp8QasRwAHH
88z/oo+dCrFmaJPmNvueuI1DxdzAzBt1+igFauEH4Orfnz6XMbG6EFJElpWb6IQD
ZvoqeKmWGeHZY6qPbalQ3S159TV20l4tpI8yWW4UgTXNBxS0f8NweltarDaZSKzE
B0U5QLRoYtC/Hm0vKENzHdLNK6SHMN29qSX7kkcDPPvUh+6s0exGrwBxpCeU73PP
d5wve+40CRTgsqVOT8fephYGv+zhINLGn+Kqdd44PcqiGyivvdB9UNWEZpHnzOc0
+26R4n1Cdep/nXo5D17Qr8GDqngq3YtkD8NfETRo/6htqrCNQGyVPRxSlfzdScP6
Nqv9l9ERVyo7Ah6h6y4kCFNG7gxFRc4I1BAnf/u8tWg50yVCFOyRDVGA7QX0B0Gd
C9sKfjIPC44fWHOVV8Hqwl+QhFy0VjQmLgvdBZyD6XkcPVqkgsEIen8ts6xR8kG0
q/VUtamFGqCu+E34m6SNZ7f83YeKALT6NiLCU501KOsO0xEYBfSkxjpdHSPbp+Mp
L1ftlVJ12NIiOgeCPP1SbfSALIlgGAD5XQJ4G7Jv6FR+4SnS+GZdJ2vkcWD/4NKX
UW8oSl343vXAMk9WocZ48ovVQIrU01LEtn71TKxB+5gJ0mE7w5ZzbNywUCNQCijk
kGXdwdrEE8DPhAzL2KVEDusy0GdwimXz0IKZjQZJOUF8ro6T4kwrOOx2tl5QGV3l
Dv5Qiw27sLmK+wac6nuNDR4TL3TpyfZyfUVtL7cjHG0iHgz4YaU2j8GItIIrkkfQ
gC0EAEdardGERI6A7t+tSwpgIL71oOYVc7ohCO3ox3ijjl4pfz7wIh1xjONJfRak
spNTVyW6d+tSMjM3JytJY6Oaj9ektEGIuXpyOs1hQYd/aDPE6NqpXO4o79Hc/MhB
DCeCtyoVuPdITn55fN42RjBWtaffr6SNsgG6OhyKs3ByBHwK7LbPdA8zPRel+MGC
TFySIiU6Acrjp+OoYRPcLsqsYJdk75xHuE8PxZZHO9HMzPDYAf9ug9sAbMkBl12o
ypka2+Ju7/jYkAiMfM1VnL0kvZVNkqh5ciMEL6tPO+c70qLmAm5T5OoPQnES0MGr
fuBdLFohykzPTmaRzFFpgOwGTDhRGWVo/CTFXtsgEtY6tn66+tgR6tiEP8qVlKR7
rQur23OEZ0pR25TO4LdV+kjWs0MUqyKWJJd+xdE9hxUwfCwe+4R9abq3HCVPSE28
HwqkwlsNoR0gRpGu/39nApmAI0FS0oo+c4kmip4y6/McwFC5r06F/Nm5dLNP/o25
IWUvDHM04s4abOx33xPDLZzR0ulR9G/bXhm0/3fvvgHaY+xOnxby8GrnyuOc7ZCv
xYn1QQdVlMesB5soAYH7Ezm248+XpHDukdQBIabwxy/17n2Q9Id729WHdyi4eS2Z
/21vd2ZIysRiDAuHXqQ6Gv/cjg5i+HD1hzWI2X5nQ0LL51gVS8ApItJjuNpmVPt5
1W+iu7sLnBf+lk/PJfQP5CEWM6Vi2rehGlue7wH/xxCoPHGcMpor30wPw023JNTG
IlelLF793yVWWUbrgcRtgugcI1y5bdOPYxsXBd4DUwMbgTbEB07FSuoVw7F3N80D
ryEeeA+O1084kZ/VxTqgdsGPMcRtw+d5G6N1oW+XB9YwR6QzUGMojbmbggBvHyZT
l6ofbNYevNBKOLV3JkpsvhOI2TFZWzsj4qIbWyYCIHQ1wl9C0QDdfTdWieGNskJ8
Wt22PkQ1//E9Ty2X2Iht84r1LwO/c6ks84bHU6y7AzZoH+YW8i4lffxZnM7gwCkt
qxzIvE6SixLpnP8Z5PasIFck4h1GRol7TyHllZsqWctvm+Sehyr2+VKb2Doq6uuM
Yrmajo51f9xWzRC8T9E/wo02dA8fGINLQVCkNftqTmoHjtxaPcrK+Mb5zyyXvfPj
naYV807RPKZQ2Of8oc0m6IM1ernxFwjUp1ZqUExnUlFzy9dkYfJcP8gldVAI6hbB
fIRp3hjkNbZrY5QaAyNEE+h9mByLwd/HheitwWJpiNUNQM+/HZg4gtwSvHkAE911
kinvlNWJhXt8bgHQZFjcursQSoBWld/Ie4/DrVwTfhqNF9UT1ZCkA9Ozmnt2z2EP
Tp1AVlCWuLe6BZD2Hdsvbae1NdHm5ozzCoExsEfnoUK5p0RMavmY+Rdx4MMnJxi7
rkdCiiNmiSUF0DTM9N1dMej2jMDVEMvRbwMeY7Mffrc9fWMs2N352x2ZZrIilwGR
jc1xj0IY8rQI1idW97jznbIG/xzKpNLNfwhfmwdQOzFzKsxGfw4UWeAQBUbG4XKI
44pmm6dDbtCRMfAYF2vTeH0Tk+5GBAveCbdJS8DJ0bshWGkMlXOnZbvw+dxRwx0C
6rb3szZUlwZGM+NiYUxXRBteFkiPqfahXmk3sNKvRP5mX+zMWnMKcmG8FnzzFIdT
lL3Fw5bJRABB1MBlqk9sDBHuK0ZZPEABa0ESIOIZnDQSsJfD/Q+I8wtlzINv3koZ
Io9yAdFB/VmQj/ub8V7EMEOKc4s6U7Xgyvx1C9RMs4b0/MI6Lwe/3oQ8aCdQyqxs
qeAlTTou96cD6Ffr+xRfOn0uG5g7LurzHcq5ARAb/PJ9QdfQpf2TH8HE31Cr4k+M
E/+A/ZR4POIsYl7dGGSBuyAypdit8lDFVzW/P0FDvBxBnk36fhIg19BlS9em1BhH
H7zWXLKWggvZRBweS718yfHj+Q32htJbr3KROzE446EUqiCLDjwRF/GuUxQDz3zY
psFXX51AUHua8/HSD4LINCuX1O8+4A/gxSYU8xrYsSsOCIqHV8EU+YgY6pWVPgox
VpboA4sFyoYSCySROPFPOcguQttZzI3JwQBPGMpraSx0zXouiIMrIyG8RAMsr8km
VooEx+jno8uKcAQQZtD4kutH2h7DynMxjjwa312SROQaixh+Gz9fOQU//ruftjXr
HNWtLv2y7w/tm55Ms3CHOm918r0xTBJJrU7POtrhOmFN3YvQlzM/8+L1jREE2/m8
wOcetZu88js+CNt8eVxE4sXA5Yob/xQPjlX6Trfz5wQkXqsZWMGI5IkvbWl5z4os
/jrsSu++hG1KsRiBHBI3eqLWRS1GOVhoGok4M4eJeEap73ozQsSfAReWYZ2lgW4r
Gomh9BN8EwbqEL45JIPnE/egWF3WJzDjq42vwYLmzbIKQdye3yMNFo0m3c8HLbJv
dVqqfD8P16xi2P+WPvdvUm/SnDdOONHcmTFHXTmwlp12tml+NRnNyljGtlk5qfkR
4Ga79QzW0D5sYoxSbwqig124nXfv9oAMwGfW2H35cfIdF3Mf7k8dPrGZdYNqXxHe
vH9vd6eE5kxsKHcqwE5V+nCCKAt7Yv1BreczdKGpIbSyVEP+awhJ8ZT3ytHzqLcO
Wf5Bb4TphLkBfe8TXSW/eY5f8U0q7cfhIIzU/3/3dLaLmLpMXFMPsJ5xKAt8uczM
nVXMKxl6vQT74xDlXTUkM9TNWBtme94NnbWr4vQJz29I+81Um+Ynv4p8jfvKNtvt
2mVJnZgPuUS7363Y3wM1eO8yZ0XOlcNwTOQIUR3FP3GBSyC0bDuh4dPOg3skpLA7
4t3q9mx/JrOYZkiCJ7V1S6nxeMOijO57Vi7EM0M1DpWZP1P5gtnGVwwie8zqls4m
CtS/UdJT5o1NNXygUeAVu6TCFBW7Oj07e6I2Q3idry1uA/kJf3xpo+vAVRFWf8cn
Iofx6AlS8fTPsrwsEaSBuKNOxMiXOHmnDfdgBbK/7wRdTwgdV72Na0HCQPdngE4m
3K+jboAMFz6z3Ntx0TBEH+mgUmjPaLijVrT5W5q5sNhfu6YwdgFZvYNjFLWSsGKv
19N74+WplfUIC1g/9DQOV44Df7C0l5uIxj4Iw4oJeCFxgcl/ct9AyFyNyWlBiYNj
RTbCXZOV04ILgNUQ/5Lgfd2HbgpNA4oarntnhJc1qWZJdAor4mAyuLuxo326S3df
+6FFBlkuJUfH7Jn5PekYnrQIy7ChHYUIuTVencN4mpr/x/6hwJr6Hl2Uu8mXV5sD
TxZXO7iN6Zvsnxfi2QC3gbO9hk8JeK2kD+a4ejJbrBrphsU64a3fQjxO2ZgcEd5U
xXAJ7nfBqJunwpH0QD8opjYs6fn7uWLQZSqTq4wZMfsRzf3Yh5VI9Lus97981Cl/
1SUL59dZzcGmvOn64vvjjk/xstXeK2Apo6P6r2RawvckXBvCfl63ZJcoOVQ/kSSK
ReBhsfvkugvURJ+O33Rdf/6sf8qE0EA84a2vDTwh6pGX/82+3kzdD6fRqzz7Mk0+
RpV8DDoJxHf9OAC26bOfELJdNLPNBtFMkDkPNcxb9rFY0hdHQ2GRYZP+9WOfq1Z1
LBXL0v3fNaLkqWtYYINJQvJq+ov/IF7t7aRFYJPY6q4gK8AzgYRfG94PSm+gi0Zx
+KdOWl0ORmJ5SWg+3nbMtD5Cz3e3zgi4uJNl6OzmohhBxeYGTc16bRNwd4pBoV29
ybAoN/PGl9xIecBz+PMuhXvL8hdagAnX5/qTLw4dRjsaMWyGDSTa257fotoktikH
+HD4aEDiWCQSTRyIslZGtYVLw/nH8Cnnies1bX5D/Lr2hwIglDmw92UyGrM9rw9q
K94uOnBcpVVarDdW+fxF+vCx32Nl5DWFehxPWkpqQX7ZjPq2Nw+8xesrAjvXJCYk
Bk7GLSKKe7SAPqulpOWmSAjTyh9FFnIj5IZRNas0onLhfdNMhsUOMGQPWCLhfTxd
P3dcLiF0xOGhi2QjwqYv4BuA1sIvLSbhz9CoaDpAnyEI9M8VWccERy/OpWCljBfk
oN9HRtSQW3BMiII2Wl/axs/qeffRFEKZjM7snyRA0Y/m4wgQJV64xuHtV9gn0Ukf
+6xim9nRa3wq7n1xFd91fv/zAzuqPHhhtQwFkl1IdlZH4Utqst0h8pFFOR/VaLSw
f6o6SxHghZefytjtlCKKK5TmAvlwZOHh8SPtNLvnT3ZMzHK4+K5Roq2GQBmOGd8y
Vk/LaZ776z97b99jPLN33KeCaM+SYVTfl1+iE1mlZQHGKP/jsfE/+Z/fvSDB/veO
i0uGY1KcSgEYncu3QQFAIIVfWNMWxCrdxHv3MkKIIpG8WDENddLN3FBdwt9wXRx2
kfaVDWvuFB5aF20x2IZUIryteLo7N0GNE8bkg76q9BBjO4TPsJnc+yChqRFIpg8w
eapYZbgOhUmdfRgaAdZxhy59og2MsIedioM6uAXSZJcOuODI6DauUb29d7OQTFhI
vOK5XLF/gIFqc8gl60/u/OcXC01GpJhakjnrk+oCESlqpv0G+CVgXPOpvjRePD//
TjzNwKbRAklLywd3M4Lt8H9wlsWlUj445DEMs1CMHR+H+yJVGLGGzM76ajszPyBk
rJHhJa4xAIZ/hn/ocKOWgs3p4124YrGV8yIElCY/dqugLd37H8yC4//3SiTKR9un
LqrMqHfdiPk3LNSYhnQcl16ygNB9obyP9DKBFu2K5ToOd92TbOYKAwW/9Dg5OMH9
3aKdWuK2PeQwTbkvySr5EUjPtGY17Fh5TnIBJtv5uIUp/SOalhn/MMJZzbCI6mN5
YgtZ7AyHuSXXBrEIp31ddvDubnaPOQ2lx3pMsUqfrDG/ny7uQiTJQKddFokYx9QB
UpZYguwg7VQMYv1UNLfcr1cVT8JoeJfdkoe2MT/6sSLUNA00MDLMw0Hxgn4uZULc
bARRUs95tcEV8YZg8DBEO89678lhypcy/UJT3qexKRZu9fUXoJsbDbR81vDvtVca
dgR5xX43X4Oqya7I97YsohDPgCxXMhv1C+TyBwDycuD+O34hYU2NOHD3ZEFm78Iu
u6cRMu5NZJQ6RGt8Gcwf3TzQZHRg44aiU7b+PPl5qONbGFITXCxZk2XQPuPvZ5Wc
ThZmTuCHqhEN/VyDttb2nsInrv+QjaDGRrzPv81m8vR4Zwx877XGvB1RkW2aEMJK
exuXJsa+uMf23zL6Xy8RuXndZ2GixuFrxG1kciKj4CvJgMnW065j34akskzGWvdE
36tv3KWyssICeKkE2gLKBdAFzSPmQwiiipXbdHiPDJPY4vGpl9C4ATF5d5/QvVXP
TkvYKC/4q29SmXUasPYqVL/DQXKdu0fOePZPfh8s9jY3CmRL8jDlfHOfIlXeAhBw
oic3yJXmdMXBtoApyqNUDf4SOxivsElPzfcGqmqYor7Flo/otf6al5F6hAZXMHEf
Qjwv4T/3on2aPZ/1/U9ygCScodBsj2krrVyuLKeOkO2Imbxg4gRePpLQE0OkpLqM
6cEWJOkOSU/0SBeN8IPLfvWRDAFz0ErjtJfOGCYVSJIyopHfPIJ2k9JCNKWSl201
yVZ7wRbqVRMOYcATccbLeXL7OdWqEVEYsG5bm1NKWjEMarYW3Tmzq5gq57d4Ah4Q
QysrINEaFTcSkfb3RNaYRRyugl2RgvMMW8F1XCVF7hwqAEG6FJliToHl5SnSzO5t
qGJNsB4J8VCNCoHwFyAOBEk8q17/c396MpsbZj0xnM3BTBe4n+1ZfQjZ58oavnT7
xvm9zQcFcciX4ZoRcYYabihY8/RXmVOfsbvDXQVrmKHvaVAXUv/pXV+63onX0Zl/
lr+dASeOzkNx9Dlj19tTWNLWbeZaOY+UfmvJCjh760MXCwVctn8idCgirGM7/yfY
Ga8S824zPMd5d81+ca+DDz/tw6MpvUCvsYnaeCk9BoWxCBVnIFSYQ8GOJ3fM8UBp
1h+a1CzUzpWCPdqUz6rZqLrLhlNnS5sXue+p4hhG8wKunhPaGuyknPIdPeZGUzM3
Jk4F7ayGAvtWJsbDhTnE7RckWz9J/QmhDzFzNtoJ2gRh5AUN8FjWS2YwIbr3MD9d
yqmyq1NRn7F9cHZd61mZUK6rH21LoteVxvs5oMKZ6dQKPhoSV2L0GMmAjFobvrOu
24nGg3HCgnUpTdBEHYrx+ThynKWm8rTOyPFwo90/Jk7QW1NrmTlcZLN0gWdzH69H
NmwNNqkQwM6iPknrI6iiu+Q4F9msrrt+/kcIAH6W91lP2SbdiD8NX3/OKzJASPBT
G5UTXo3/IoagWKITixrjUln2kiOhgmPxuCdQLJcIyRkeY3gxJvsA23m5HpKrQzgm
RhBXxdjaDCiIi0NbCDMxqhjPGijX4w7ra1GHI1qhx7NapRdk5ucrbo2hRfXpLXlB
tQZDJ2mgucEiw+yBoGshcI1RN+qn+XBufv3lUebvlj0Xrj6OaUkFbtsHnt2khZbM
QgoYmBi8dAvS6vpzy/VX9vfDXrgMLuwV3BLHu2FtVbPn9uRqEjBHQt6tiYlPwm7p
0SYP/91WGXzUgv9drYz3eo38ZrmPTKxYUCzaLx/18aU9+GKXj9ZGmvfjJeTPwQB0
o7zhDJJcrceUXFhOg2GjpKFSuY4s4mKMZh+Zh8kjl7yUBWUJvCcU6phKbWgq2l24
YHkhakn2rwDyl5uUPHafRoPpl7MFjlG/jLimBRCWRD2dZnZ0GNoh1/F4BWzsZE7b
vpm81n4Y8IaP+UJN1pRm0gmmCL4BjGIzUpcJMNTqzIAAVbPS84v+O0e2DAjWU7+O
h8r6beKLQdsRc8mSG4OZ7marvRXEKbXRkO99JcIFO5KLaX2VGxOwLyBbrhx3/oao
FEqeYPlulq1Pw2dzC3vsjx1NIJebVx7XfRlojbHncAaTlSk+zFbrliBUvj/w6gMw
9j9IujhDV772Zvtv0yMiBv+DfqTBRmufQ1PokVL6YMhx8FJFFLoHr6yXmg6hnqh2
jZKKODyO7llLbsI18OmjxbhJ7lkCJdUjlvJXlokqe6np3Jfa/HfeZJOfHNwyOpGL
TDXx6c1+YMIQ+31FDj42jrMR/0GA17K/mgOailBHW/BZNCGAaZA56C7liD/2k1Rc
0E+/yJ5LDrPm+BG1YEOSR2U7GkPsuug3hHVnq0jW1TKBS9Xcog3BKrYZk5x7yHeH
P2h9YF5ZDidF7PnAAEw4Zwh6WOjD6VMwBlIZs6ckxRhtYcQJliwf90Q2/nby0LgH
k5oyUZPO3hMEkOCGi+epqqm7lI9laci9fVp983418iuJulqY0f1kq+2sKLLx/lXi
0DUjQLJeX3L72QOBtUlG/z/6G1gGiNkT5Xahgvc1QHB7OF1FdUQJ+KIlLw5r4tmC
mH60XUD1JguJLIQsr5RLwv7nADIWzNJlTOs1cmKhtRx7nSDIftzVAxNkw+sn1Gmd
A8AvbSwDMp2M2gx+n3zsOG37mWEw0Tc+3fToQUrs2we2Il30N06aegQjfGtVNOG2
vLUArslHxWAczrepWS5Ii948Qx4UjB37HuuZP7Qfsm831dgKo2St9X15KYa1k05s
hX42xsp3tCwe5/L6z3Ab7jcQ9iHd6cNJM+A/1SP4Q7mleRgf/OrVutIwBIFlrbXv
+Le6w6aZaoi1Bw9FXnsvkgjII4018KL/2NklYj8hFhNOIKISWv76LJZmpzjRnXbP
YDnrv8b97VEdaq7CHoUawh7rmsw3E8D9jAzo3rCkkN8xnDrqDmp8nbTYO8kE0hTc
tVEQLODQmX3yKdAuy+zELX07jWoFReIgiUV/uQvRRCouZwyhw5HfJcdszhWxLmfr
+tuIroU5IImqBoT82LqOZ15HSty+1TqYQ1rrDaM0OCeMOoomkDxapZGe6q/3iw+2
N2CKG/sFCRVNPcRfOTtfzOdi6vnO0fxADql19sL3hWZZm7+QqkALMXltWIfr/R6L
GkDnUXD/lq6T4RI8YqJp6Dcwlci7DiGO+M25hGVsJb35z1VC4YhkuzDP+vn7AHyl
QVXrpW9V0Ke4BM2MGfPQIjec7tuwou0qoj4krE+q5/zQ81VyMtb2dT53Q/7VgE8D
55fnPa8fdS2h+2giStSDRKqhNgDKQ1MODiXmW+wKpfSJi0atCq9JmkxZhq59MxsX
3UpFEyeELDRUpv2sRmJivQbWzwiEhM5hqewEsHVzsboHqEqU2+2rhu6kK0Y6YW97
YEMNOdtOR/Z8OespVfUUAf6PuYOxD0F3jOS9Xln88wgY5K/E+MytPk0ZCMSlCHQy
O2f/PDtRs2Q9DzjxfR7BHadvtuxNwCUnwewUTbNy5vbcC5FPHB+TlGGEzd24sh9T
luvV9Ikkr9uUc0fPEokheOF7OD+eKfhWS4FvEBqypWH2mgNczd6BICFR+kb5A3Ao
7q6Al5dRzjbn7p1ZrbsFZky4C6qpL1aB32l5G9zv6wgDi46ZIwsFqSJFHXygNLFN
drnszbK98xTZJKL5xy8IRcqVh+AUMS/4KPQfwgaEGa59Vy+EeoV74hL/KtpFuYpu
Qfb1pAatVrwCI30LhwMRxB5SC7TYlFK2YmFkp9YXlMh0LefEkCXMSJhjn+zJWKuf
QXJfBD3l48/Jsj0XmLINNtZbewH4q8YWgV7G3leNkwRDKhFI7G43Cz4GwmoCK8+c
AP0MpN5N6pqgYWe0TX4m4YzPQwDO8WUV+ONwiFp+WYdEnSTGIp8YvOsGj/4ygpZv
aBLciz+bMQ5EMRDM1zaKi5x+6fx/IWlGDDezeAxzombVbGeg/sf3FZjiHy3l7vZl
iNCq5QZFpBEBEMw9x/18klku4U98aCaEP8Q3OOqGIHb6pe18Aj6EUpzyfTDqvq3T
x5FKqRy/FR11FvOxYtsJp3zjN6Y+1ZMF+uJM48M5LYml11wP+aBkZC8XDp3yMTNY
4xl1rOl6JXg3OiUTUtpxzLP8eUy5rkNua6Aisl5q/SFxqKLYlgy/Juyk16lABQPn
oKvyHZPREJqM4fOBD2zN0smNPdGwVDeuNvuB7CiZG4QtBHM2WvK//gc4fpt6zJct
t/nhha52hUMfW1EfPRUqLpa2Dz5F9c4kI2rGfz8Y/HaRvLfpQQzovLJ2L+9dIVAd
08FjlFUZjSb7xNS0/qjpqxAVSg5UCG68WFX+G0ixcXd0tD1lAsWhNOA0gBybogxW
HyjzF+S6Uvn1CHJayS9xhEZHn5uGytLzthtzgN7r2YlTvBxiV5kNZhHvI0rTRVNy
VK449Ew6prvG85wM3HJZMbLdpOpkbBFL+fsLtxtJdQ9V4LhY9pFR9PSA6ZERfgKn
HvtV6h9eQCvw+irPh1Cdq+AdagvRbHu1mvTBolBhDdMnJ4GIRmtDdsxZuVB000H1
aaS1jODuyIGpX8rrsPdrgbzNH5roiVsp6gY9tLS7GjDNvBcINM9hI+1Y3Blrxen+
RGWj5bd+dG5/99hbRKr09V6RzIhnRU9ffoNYq0Aiqgk4Y4gHl92yR5W0n3p1H0vm
ZHkz2WeaR3tmw8LLjnQaDu0JcbbvUdNcObjIOmGyvZQHoEppzKJz7lODMeTBYxe5
JXb0Pma1bQ+Y+q6iz/ELGBgXtADqRn0sDdt6h6+PBJkJVPvemO8P6ErdiEX0oewc
zfm8x2cR/X6esf2cly9dwfaYW8wt+O4lAQBEg/Mt2J4raJ5ALlAUoQ/E7xeXQeLH
Mz+T3+t3mU2hdFLqQyOnb4y8060kUTShdajpaL5pAltXgoxjFCZGW2oxBckxMsxI
0EkrK9rPD3xLDcjfeUWdoU9SpWy3I5jjT/OtMBUnjajDz4hlXJqjAYOsZ7nx5UGj
ELusjH6Tz17HshVUDRlbjIAx6zwHU5mDPST2kCC71bKEGD3iPPaJPMgObXAgT+lu
+8EVFa8UJjLuYM63lneFeL2nrgoz0Eqq3j2sakY4Ik+QYhjmB2a92i3aqI0NUikf
KGbC1x+fF3weoUFKC9d1rKecqvjGxf4y52lVgK+0WQ9fennk+UAW2r9f1sgG8Qer
GR3fA6hcKGaD+/KV8SJ+my0H3ooZPfLWOeBrc+X8crCSF13ptqHssYnM2j04tVQC
tPmM7A82wz6vHHefXi5nvZdDar9qOrKUESA+HhVYdHsd377guyYMQtaNRbZ3Zuxz
Dpw4NXD4KVSt3H76e5dd6cjMEpgTG4rJLw6ZYo4Zb80f8vwsJQkouWzeVjgPh0kx
9T66M7S+wIdy0LBsqzjEkrLJ4fkumNjjOtgdBnAlis0UJXajTRk5FZpP0LmK0nfR
8BJPD7E9obnbu+8dEGRjAxyxKtK7CBsJq9aFlLrEOeI1kFXNFpE88GNUXhencpLk
ILx9Zk/UoB4/pg+3dxxzcXXLp+ascW3nHr9yKn72Zue+roNzaxibSeqa06EgsqFz
y1qbm765PX9boYG7XGWUhTQYKLskJAee77GcPkqUg3R/VNi34cHrZNvcFNKe0eJK
GFxzj0cdztdLMPHISP5Ocoxgsg+NLCrwdlCnUbOnvhf495ze8d7OUdUwZ8kxdiIF
h64aBV5lZ2natdmY2a5r+8h9D/F9L1LTH3IW3dDadOFZ4urpKPy3XcXh1GjH7qmm
obupw5X91vouUbGgYV9RjGTeu84wjIsYig9Li3twRtfvydQ1qB8qur3wkKPaUz4m
q7m3y6mJSzabcrHas9yTLvEby0oRqzrpgU71yRgrQN4elcXXBhbZ8V3GVzVFlgYU
qRzSpnreSPte59P8CmpGJgaszeHMhcoNxXxcZogtexN+38khav1IjSzHtH4VuVoI
e/T1I5KrbNjucADu3VzNW9wIWOw2hJhTmtvM2jHVBa1i7IN0xYK1uOWnhxUPm+Mc
qAQErLOfalu6M2LaabU02ECZal+teqG1UGdkYk+jnrXdA1LUfkEfF0ikY3++DNLk
t+gMdAVB1DYt/Z10HU9DyhXJvOnaqmeVHm7zFgdNBh7jx2EoqBcLqZnbdrIzllTx
MDAdygnZRvGQK8A/FlFfV1/oIDV5WBmYTz/6bGZ/MSdU9cBswhJeNGgI+YLKMmeP
Mxhx9xLHFfErh8KsrEzXdO4y1NCAGqAbM0Y4O/HhRbmYHReUUOwPbgGA971HtjmA
gY5McIWGvCQulRHjHmkQaaITQUgFidaiWL2t/ONMqiPbk/TuLNzCeelL1zTjQNzS
kbaeD7TzXoaZSBfx2BOO1XYUKjlEToHqUwJbNNPuS5gMb4tvJgJ/J6Bj3knYflK6
oCwPBlwqlAGSiVzVUhz6+2UDFvD/WFjO/Yv44O6uEMPxcIawQyzTeMTnDoKIox1n
i6m61FGo+6BbEwpQkuQET9AmLa+b4+LblZXbWjAOgWvskbUuxdHQqDNBogG4bYCb
F5ySSWYb3jHa1jBMZMIld7djl7bspdrZxyxsL2/YL9VRTs2iUXfbC+wdY4P0fTBw
7YXDWqNM5+ob37ekZ2ZbhtumOtGnqH3lm774d26oa7aMjp0oBjGVdUmTmCnX94Bt
dVaTsH0di+VJr36c1weT1cCuWwLrVfeRKpopAiRJRdg69s0FgeOPTgrb1OUUzf7F
hq9VckY0RPKCj9o3NruSLBv76955drGpt4Ozd52UZ8AdMCnC8AI+oRzgNzG6l/bO
ugVmBgAkCbVIxtoROf+eyOrcA9mSjr835VzHtBa9pseJCguiklDwE4e9KHryBKJ7
7Vjs4f/sF6feiUi2kOpXbPS547wDRk1Lk9PxvqCcJBB8zOsAdY4bnwk118IkH2NS
rYeLLMKfP0Ij4lugHKk+Iq2xCfHIeEJQHQaKIG+oDPrNknHyPf5+xEFHw9mnfx3F
9SaNUZ84ZSsxr0y14oRN89MvwiUHLppeS3N/eclKnpY66rPALR3HAC+X2kX3HxUY
cBb45COyWmCXji83th7VD8F5vxbfQRRVW2lHPvF3epXx66g1aRZaB67jX0/4E2gd
SYmn0ffAcTIyrqJviNa7ECNT1TyFddtDUT/u0XeEB5BwGrR5ud4Cpx4URqrbDS4T
6WgmI5BkB64k7DLAQ7YB1sx8VE9ro18m8D/F1iCo4oBs+E8ifKh0tJ0jYiRo3XSn
58CdrqVgsn09YYxX4KPfrMph6WF5iS69n28xZFG8ziMklTg3lm6LvqmeYCXC/Ini
a6gDCB5cIGaVuS8huzFU0yTfhEY47X7axxSXjBDXY7avWDOU/fBNrrDgKK7unXec
beMKjrHQFq5yeqxok93LLTjU/roCXZuL573YcV+bZ2BMrm9O+3DU9hjyI1q02hRw
6InqZheGOMasCgWFxiYNmS9xjSELqZ/2N84cHCaZb52i2iUPaaqD3Uvwfrb9Iafw
+h+Z2NUF9R5lXZYyK1wEHUwEVsJLkRsFXCO4tOaGfr0YkoI9kix/IrNbqJ/naWSu
CHxKHGtd0pAsVhrSRQ1uFwRKx+ETvR9Z37IZzUPNJxoEjpr0ofATbDBD0s1y3Joo
VBh6MeUf+00lGPFlpZAp7R3rt3gSnqre4jPAe2BqwXoYQz9iaP48tpvoKYLjKuM1
abRoT0+Lqc0jmBjiJlfgSpueufX74jfdtGfdTIoRytxv4Zx8unIqrykHbfsCTCVq
vqcQ1v4Fcx0oCnw2MH8wuIQx//kZNrGPrKNGrIYVexxcAtCNzdrIKvK6IjVVfD1F
qmI/0KRJJgUId9m0Fr3VoM0FNZnBtxbZxO/OZw6f5Hh/hU0GiL65eOQdYnol5zJv
O7ZPF6jaZkqcHFJ77LyOWb45u5WwjmRKIC9ytBpyEElqV+PydJb9B7tN3z4xskWR
ceIiBpletrxUO67FJGH/cild9Z9YVOII1u3Y3s8T8F2wWHGEe/0sKnu4+AQ01YS2
HEeT56uyFEbRxGmdm+S9jm5pFezrlpftfZBf0Shbg1n35LuVqKmTFMlxoSM74IQe
gSaw+EdWSwFIpmGs+Xo8DhCWIqu6HiVkINVbrKvdN4jzJhJJOavQiyi6ZzGtbpF1
TIzXYPuSQyWhIM3UcCPy4j38vgWGDwzsptiz0SR2Ei+elc2ribFMaTNe/IHuuCdA
q3JMMZdP8ZZM3zzhHTA6Pu+vYQf0jsiDEYxJZOGrDEHdUWyAwZvp+ZEaEzhtG4ZB
D566K4eZexeIyN/Iv41tGVCYm4Ez6770jzDchXDswjExgab17EAVrkrruxiqAQY6
TyBZbUy6V5KJBjVs1ZwFD0bIn8tpQKdulrhz3jIqwo769BRp+FCvj73whKvpwFCS
tlrS/hNxtZfPjS82PAISogxzSuzl1QqxRUDFgqEFRfIcAxaMil7zG+2Qb5g/7u7v
BxxJWxvj5jr3D6GfA1CFocSVfXeLTvOEqyTDcAhEQHTUIdqFCXBGVrFGZ/iT63+O
NHaWaPxV0BEZc+UOjtjoCIQ1lWFpLpgjpZfvSAtbbyiyrPwYRaOoog7N3AS+uf1a
EHrbMW6/PRonY5Abdr0YuOwqSH162HeMinM7ayQrAVnKNUBStJRXxq3r0HtrTfCs
yzj2cuL91JRns2lWI2PK5kMpO/QTqaBRM8xoz61eDo7BWhbYqHl8lpGWbIjJSrJp
bRewrHJvoVAQCjb5ibDKqyfE7pTHZKRDdIYarqTTFTjAal9aDlPjmz82CK83iDPn
DP6Eey/XBxpeO9d2WUy+kSOdt42yoySeUDhq5X02Yh6XY4BaNBjBUf91+oZPDwC7
aMdGEo63mWeUOOcbGglx5KpoMjv/lkmfsBTDpartv3zl7okW7eNsadRqxdUPhU2J
tMUTaI0+VGY7342iA7X3NCtHLl/pd6HIaK8Wzgy/5Q41S9BZGEY7iMGUo11865Ye
VooGRtRj3CTGyKSEi+qDBHVHAxwvs0xS+WeItZhSgtgSAdLon1SQNzvvgnvksjSi
v5uUh5vnY9OnUzfSF3v98AR4faBSu1IUYTetn0Vo84tzBs+OrenrTBj0qb5PDDUg
KEeXNcJ7W0zVOPvAE7X6JNfKt6G/D0EUXOf7LYp5pX/5AwM/P2eklU2T/l7QcaI6
N1IMl4DjwnzmBUgHyia8nsQ1v1kmP5meN4aXzCY7lbMM5IhFa1B2Hd+JOc/t9489
5h/LM7ACAAL11qNrIqv8gdUCLYAK7s6us+alXqg1j8UHQsFTcIM9PJ8P3nNLw1Fl
QDq+4OOg38jtFuyjGf9QLNwDEFUShdNoJXMArjRjwoiR02CY4kBAp34qlOk1uSOx
Fcc4poI6OggGh5Nh8ZnXmXsy/j9MuZvr8D9jdbY3550cQc85PZeelO1UPzVv3gQj
si/OIm+n1BR4axQ3VLr2gTeN/9Nu4Ke32Nd/rLAriKOXN1LsHdiJOXN12M5pvGzl
nPczWDy9QPNFllCiJS3JVjei20KFcTQb8AiU23K7+cnN98zuqFY9cxExZao3i+lw
G1yeV9QGjBHNoKdPR3bMftFUzwPpvP4b73eaCQxO6geZdgEhnI5UiflnMm3/xdG0
nI+mB9KmvhZ5+0ezgadLk2tALB5oAH2hW9M6K1J086A4McAbUfTn1lN/vPPUC49T
PFc17U+ma1L2ORDUHEyanKeA6yDQOX9aZHAxevFJ4qIs1NX5H+DKq8Ct0A8arJ7q
33T067DPUT3zGiDqyor/3v+4vSyFvfdzRb9UQpRA9LSqU4EYB4h8p2fQTUHQacjX
qoAyjTj5kr8nmXwaWJUXEG7MoOVW4rd/Fda9846BaKFD6fIXSSCukQiyOlgbQJ3A
fF47L0sDzLOv0Yr5G8FmCc1qbMVyhLFyLxJMD3EOtSyLhKYUEsjrSwZK8B4ToDvK
xixuMlsXPhhB+SvSWBnYz0ei+SjB9p1nmnuscpFtplzt1VgFFEhqQtUt0SlG43hb
5dTG01lPxKEzbGB0yqVnq0rcsbCCI1wWgODgEU7rbOm4UvJZ3A0zI752XR2I49Pr
uX2nTpW+o8NC4o3Is8HOFLuvqya9PAGzFIO8aZ3aLMWisttq/B0GXLf08tQ31eUh
Slv1Ok6vZJsP1eNakhbcqNYsImCzFEnHuDAuv+Z1/FvgFdLA5T6gLWg7A0qSplOq
rXqaVke+qc+Q4upRcZNGqile9RWWfENq4/efCnq62qgSCAAgcnHeXF6F5s1ZNjkd
3SQGxgaJST1v9WJb1/pEP0GqK49lcqXft6v6zBwwlgwMogdsip4A+zl0g1FFsgPt
HD6VVd5tp1fsguYDcipB8CK+1FWGJir03AKF2Mwev68d6ZdT4KOfr3k4f/YUtGY2
vcMnnq8HCMy2GXPYNwtvSWvXN2hXLXCJadx/ghjIZ4BJ/lkNBwXznjNy3+G97Glj
V69tw2Ee1fQ7FHmhOrcvxBxEMzIfwuFaxcznjylSjYoN+ApcrOIKRTNwPxUpABKv
tpbsSkaWjO5IRSX4V34Gz0Lclh0HeB633RUYUq4oWRvQhb90xtPmAbbth/dtJPsD
DG6BKiBKc2OrduqFC5ZGkhsHZ4sGPa0lJS6WOU27dyntpACgJ9BIkzrfBgMxw0yB
1SRzRFSxlOC+gRqZSBbOgniQoffpH6VSghngmlzsEFGItTRzDP1vLb9YlW8KZ3Y0
1mn6gCopVitGszw65diAW6mLiJYwVPVOTItSZcgJU7bBOqrL573x3r0Z/FMQxxl8
4oDcSbj+nD++P/EvwG+0Uo3FbOixCvG8E7OtTHVGBA3SwQKZfOTJzIQRj5MSDdiD
qkaukwlFiQUu1CTUKHPO7D1zwA2kCBqxltMMoJ5h1yV4bmluAJ+uLDj2bB69WMUx
NENoh//BbtD0QpPhfOy+m0vsOnG2Xjmp2UwKImZeYwSmOBrQxrsMNBzPqH2x+A7z
jg9DMr3iZJU29qQZjeM1pgV1gaYoeLoTMec9ZgRM61aVFf6xJ+M3Gff51tXm9Pt7
bAce/3HXW2GFFgR8Qeoei44UYTBEMqyeNBqOn/4UC+ZuYymoFD9G8NTy3IlSGi8N
fcKodf2w9Hp+rw7FvyvVJNbvZGl8oeKw1pxUgGxUUV3E57IlGY88yZNdIXLn7Q0C
xRodH8t6J5jW2m6mBFuASr0tiuW//ndKuvKL+rR4/wnjy9FBafAeH2Ar4HUXvnFQ
LK48xnGBLa9BwU/4DcCJ5F6izE9O7T7mSWEVJjtAKlkODAHexq7Y+oDXVR2MG3hG
iYlMjk+LuUMJ49nRVWoG/lJGVfsEoClKDPh9F+xJ4dD0rV1LsYCsRoEYDI7pT6bM
cbNvrdKZfdsnwGleSHf/vhFfUjwqJnRotzzkWC7JnH3PP7q2QiZyJsWWvg2dzQhx
aIEjtHU3AjTK7Gn677mZac0g9xsFc20kKI0MpkiPK2zmh9jgzWQXVI8GJzKI4Xt9
m0W6Kxq0089TuLYAxgH61q2BtrfBlmuUBkOOmOtviP/e5kfE/rOyxgtu+5bH6scP
9wyrCiwZREmoVKqv14O61eEmhW5scqWR3rj3zYGirHkNtxnHv8OLnRbBOJxo0abD
aR5C+xMMkdtqI5KTbzpGeNrX5bKNnhzFb9gMnD49PLSajGCCzO2ghZNr5viCT7wO
pTVLSou79vOKlpcwkOTAFjhgzf1RQYFuerGzwEgIbxrfkDlb+3e2ShyGsY8foIOi
YSS4LoOwxcBAjKu1qTP+q0z1p441bqA264A/+98HRXjGWHHQMtWBd+qACEfHOmlE
Of+RiC00fxSF+25iuQkaHYwoP4SQriafiNBD+ZLSx/gpCKEGWydvBa/8nfF8Rcaw
Ox9sUtWIzDNp16dg2RZh7UGTjRhGNIoOT73Pd2u654mDWDtkMgZLhARvGy7xz8da
P9c9eSZDit1N570tP4QwiK30SNlx1bQ8cRIDqCt6jead4l6nGKVFBg6AKiVpgDyn
d3F19D3m3VuzLoD7HMvAsgkhRf3BCpsVi2+U2sjA1bOcPSvLJI1oA4UngVQ70rbu
Pa95n5Mw5vl7SFE295KiqCqZii0h9Xi/Om8u/4hfDsh/MNRZcEF2qyxIaesS5SqI
HYuWyKbvsZAI0xxtk1/scbr60BB1cn+Iuu/RA59SDOe//UMuiXjrNLZKUv1yw5Nf
VWUg4ODMbQ3IP3EHF6UwBAuOYJQRRBUuCJTjOrdvgx9Es3tYEnXbnLla7UORuKED
nXlWoXJ9t2jD27ZATkj7El+QuaGBO42DhWlAkZgrSL8mqBoQdoeDKm+cvMUZsLtr
6nkyFkhi1JUcnvcaNu2x83MkIYNWep1WmgC7r9/yyh5P5C305eB5aEUqeXuYSmw1
ph1kkX3/z0S85O7K2101lhiR9kt6a4nk4sW/hLtr0eKcbwQf81pYyTrVPUEgFKRd
u0Qky2iOzTctdKhWcyus0Mao3qnr8DCfaR5L+Yh1UBtgyJ1zrVy9FtcRQ4OGB+Z3

//pragma protect end_data_block
//pragma protect digest_block
0wMPYY95W9tMWM+usmw2jIBW/mo=
//pragma protect end_digest_block
//pragma protect end_protected
