`ifdef RTL
`define CYCLE_TIME 4.5
`endif
`ifdef GATE
`define CYCLE_TIME 4.5
`endif


`ifdef FUNC
`define PAT_NUM 200
`endif
`ifdef PERF
`define PAT_NUM 100
`endif

`include "../00_TESTBED/MEM_MAP_define.v"
`include "../00_TESTBED/pseudo_DRAM1.v"
`include "../00_TESTBED/pseudo_DRAM_read.v"

module PATTERN #(parameter ID_WIDTH=4, DATA_WIDTH=32, ADDR_WIDTH=32, DRAM_NUMBER=2, WRIT_NUMBER=1)(
        
				clk,	
			  rst_n,	
	
			  PADDR,
			 PRDATA,
			  PSELx, 
			PENABLE, 
			 PWRITE, 
			 PREADY,  
	

         awid_s_inf,
       awaddr_s_inf,
       awsize_s_inf,
      awburst_s_inf,
        awlen_s_inf,
      awvalid_s_inf,
      awready_s_inf,
                    
        wdata_s_inf,
        wlast_s_inf,
       wvalid_s_inf,
       wready_s_inf,
                    
          bid_s_inf,
        bresp_s_inf,
       bvalid_s_inf,
       bready_s_inf,
                    
         arid_s_inf,
       araddr_s_inf,
        arlen_s_inf,
       arsize_s_inf,
      arburst_s_inf,
      arvalid_s_inf,
                    
      arready_s_inf, 
          rid_s_inf,
        rdata_s_inf,
        rresp_s_inf,
        rlast_s_inf,
       rvalid_s_inf,
       rready_s_inf 
             );




//Connection wires
output reg			  clk,rst_n;
        
// -----------------------------
// APB channel 
//output wire [ADDR_WIDTH-1:0] 	   PADDR;
//input wire [DATA_WIDTH-1:0]  	  PRDATA;
//output wire			    	  	   PSELx;
//output wire		                 PENABLE;
//output wire 		              PWRITE;
//input wire 			              PREADY;
// -----------------------------
// APB channel 
output reg [ADDR_WIDTH-1:0] 	   PADDR;
input wire [DATA_WIDTH-1:0]  	  PRDATA;
output reg			    	  	   PSELx;
output reg		                 PENABLE;
output reg 		              PWRITE;
input wire 			              PREADY;




// axi write address channel 
input wire [WRIT_NUMBER * ID_WIDTH-1:0]        awid_s_inf;
input wire [WRIT_NUMBER * ADDR_WIDTH-1:0]    awaddr_s_inf;
input wire [WRIT_NUMBER * 3 -1:0]            awsize_s_inf;
input wire [WRIT_NUMBER * 2 -1:0]           awburst_s_inf;
input wire [WRIT_NUMBER * 4 -1:0]             awlen_s_inf;
input wire [WRIT_NUMBER-1:0]                awvalid_s_inf;
output wire [WRIT_NUMBER-1:0]               awready_s_inf;
// axi write data channel 
input wire [WRIT_NUMBER * DATA_WIDTH-1:0]     wdata_s_inf;
input wire [WRIT_NUMBER-1:0]                  wlast_s_inf;
input wire [WRIT_NUMBER-1:0]                 wvalid_s_inf;
output wire [WRIT_NUMBER-1:0]                wready_s_inf;
// axi write response channel
output wire [WRIT_NUMBER * ID_WIDTH-1:0]         bid_s_inf;
output wire [WRIT_NUMBER * 2 -1:0]             bresp_s_inf;
output wire [WRIT_NUMBER-1:0]             	  bvalid_s_inf;
input wire [WRIT_NUMBER-1:0]                  bready_s_inf;
// -----------------------------
// axi read address channel 
input wire [DRAM_NUMBER * ID_WIDTH-1:0]       arid_s_inf;
input wire [DRAM_NUMBER * ADDR_WIDTH-1:0]   araddr_s_inf;
input wire [DRAM_NUMBER * 4 -1:0]            arlen_s_inf;
input wire [DRAM_NUMBER * 3 -1:0]           arsize_s_inf;
input wire [DRAM_NUMBER * 2 -1:0]          arburst_s_inf;
input wire [DRAM_NUMBER-1:0]               arvalid_s_inf;
output wire [DRAM_NUMBER-1:0]              arready_s_inf;
// -----------------------------
// axi read data channel 
output wire [DRAM_NUMBER * ID_WIDTH-1:0]         rid_s_inf;
output wire [DRAM_NUMBER * DATA_WIDTH-1:0]     rdata_s_inf;
output wire [DRAM_NUMBER * 2 -1:0]             rresp_s_inf;
output wire [DRAM_NUMBER-1:0]                  rlast_s_inf;
output wire [DRAM_NUMBER-1:0]                 rvalid_s_inf;
input wire [DRAM_NUMBER-1:0]                  rready_s_inf;
// -----------------------------







//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Tdl91U/4LkOdJGo7eLIkfICNHD4aDqzkPNPsdwmbqgPbhLNXTGjhiT/lCfazEG5d
/J0VoU1SmfaivBOeiDR2v4m4TT1IcuoVLq8/BdxuW9mqtNQDllKwv0UzoBAwhcIN
Go8yDcub9FJnc4KYkqYzpbu65NjAN6uGDWtVqgIcuc/bK+CHFQhJvA==
//pragma protect end_key_block
//pragma protect digest_block
Fxo6vFugXddiFBbPIVGCZ1yPN4Y=
//pragma protect end_digest_block
//pragma protect data_block
vPpshDXr1/aGvH0PVmrZ77wTSZdgPWaNCkgk9Mq9+Ogj2I7LqahbousbK1KA4cnr
5OV1J2Cx+OpwdhIrdrLSwY1imxSNkP9jwhBC7QCD+dD/0sFaiST8SVV2vKkYhMh+
9XAxFvPvHJqckGzRPJyNK1f+Xg3F66+OgkzyYBJ6J7yLwtvBuyFt+ElJ/QKHpvjQ
ZgnX6OowPU/DfUZ5R+J29tnfx0Uk1BTrcP2Ztsj0Oe1wVmRaBx6gA0AQooCU+jTY
WUBDsTygtwPzXlBDBuI0WcmOlGOO4KZOQq2CZW4ljp1m4E7xcAJVR4g+59eLqv7y
l7jci4GfbRboEwAid3QImk2N+vISB2Vf7ftTPjefocC3lIg5y12LH6xP8P/XT3/+
1733QoXs6o9puawjHUC4HN2YCPM1XT75EiMQlxlOKkdlTY6JL6ymWI+oEsyizs4M
kut4LRw2LI91IrK6kaKdqsBZuOZCRGKjCBgR1RuGwGQu4j3O4CPOqeOCpwGblZSP
GnyVwpkEBBrtUIhkiLDIKvZ4Za7IGkNTVlCl+LbxbgNrcWkpep1IsktdlWqgzB4x
UezHMlDCngBBdatPkS30gcno9xb06q9Fnqrz71uW4s4XfQI+IXu2rsCHA3x2isIE
TTij7kim1R0FSpU+KwL9HOgqP5Bx0pSgqko+o6C1jhb5oHPSCqvWcdyBM5pG3JpB
L9pzHcjgdMuXYET7BLJNcA+CGQnZeYd2lvBPhYwaV3L376tnUF+u53bLz/FCdk9N
K7vIljsQGloenGfbGjz1XrzNKsWKxE39q7W8O0dEis3+piM8YvcIXl+6veLA802L
raez8w55vgUouY5Sw8IpbUNImx6GYVTNDynXpFuvUtsI6blH4JNgMjOJ5OR064Hv
ujbfzulgwYWwdD97g8S8yuj//1cBhhUkM4/D8WpwP7iDx+N2IVHZysGIKzL+4bt/
7AsEjF0yL/0wshCD5JK3pZadkRb3e/83k9hK5FNNrtAvQaSmknbkaTnUbaHzCR/7
oU86rHLHNFHWVHTPEGKWjOm8t7PVr9ufxX0ayZLyNo+Nrmi4QF4xGM8GaXWGBjX1
0inV3pFB1+appuOwSsaEUGSdZzjGpbERLuhTdWgk/jpfbPhROnD7wmIcsH5yynIL
JWl0xJDbKQSXAJfBBxUq0h4+uoKKGQ7Kte6kV1dU8FYiQdYYUy9taTbRzijPbYNN
xt/vInhbpBpT7qPNpfF6Pnh+7URrAuOwtftFtD+NawpTxAqJ2s+PK1IyRydQTXoI
Y9uf+5wYFkFatec/h3VM/9dVNvYqis3QF7v9NiVSYu52ytUCXFoN/M/47au8LmNn
fz1BzxD5S3KYJCtMemtdF4pvwTQGw4WmcUQH9ITlFSB17gCzcAaiXkOp3H0yUOQq
Wfwxla1l5HxvKTpJTtiOFxLzMGaABjB+Gy6+QVt5UztOeYZhIUL6e3WhsYz8Cn3H
sSSmIlKuvjDoWIblcy40qGcFwsPmvv26sHff4IFe/gIC5L/cNOPWujymT9egZbI6
iyJ3oDiFKYxXN0HN3tWu49vFbmz5wPl9jZIFM+31c1CwPy+wSZQvww1CoALbaKKM
3vvMjkYk74UwzV5xaj2lB7OYmf+Vl2cXSmhOTSt1kUyTBtLwgWOcwOeS8OL6AxIf
zgduPTdxmajxF2FsLfyk888ZURg/t4PnYbxSjeaHL3ndthPHtKHnY+wKzJIVBWtl
fFy6xIx2kkMo+fJB9c8Eqd50QTrq0jqc3WBqo3XD7l+cd84mY8Noo3RzdPFk8XLk
/Zw1FYbHwRcfUQl4yzgjMcW7jXX5EMbh+jw/YAk+1Hxmu+L7LOEzRvaStPAsKlZk
kf2JgTTnk2fg8fIFCG/TtVFv7NQecKgLv3JGTLPtscQBy2TFmikgK7j1Z5kImVdn
E4KDubInnVaM+mctFW/gZHIUDg9H9+CFV/YKbXvJT9jK2a9IC5dxzeqzCsJ7jz52
M+xe673FQ+TAbBTm8tbTghOMHgqx35tEjsXPoxrkF42MFp6aI/jRVsugPclvBfnY
TwDbTqNj4VCzxkwdtY0Kry5NKvcxTO62WKxSgCZh4ikN5jDpYbboZCzMjMd1/jK2
uq2xeDsUaPgAK3TGl7LMhTOm61l1XfS+TN3ndMhT++jMptGhRtLiOj2i6OaXcgaA
R21q9INzlSGVBoZw2rLB/xvNXKo1pNss6UNN59p7ir76xaHI0/b4Dl1PtTJ0WOvf
UBo2X3n7KaIUiysOLrdbTLjGEMTQnHybnB4FeeqBeiF/ftWaKooMCX5sNHs0QByt
axNYSVYNZDIofBBH+yz2B/klnt8o2Gd+pRYoiMFU5zt4SjXwWR06FgQbceZ+dRyP
xIAviFwjuqxaH8yyX5iUi3UWRMh5fIvuW8GiVJaQx4K6irG25Rdhv8dhOSZ2ffy7
22E02XZHKfy6NEB05Vy5If8lIRmFeqaLvcxYpmO4kR/JKMl7HFeBGb5RDyGvKM1I
ZLdldv87xx0banYKMFShonhwwCFFCTjucfk7Pu5OAbgjjbRSyJ/MKi4o506Xplg4
v2SxK+ue4OhfZngZhwXdZxcN8tqnvzDC6STK3cVPncfuozxeMOehWYSYgY6prPKb
ENBrqmEDCeQ/NT8AVSNcjSUgyUnPIF/girkeZqWboBHQ+IuzTgxcr440dAB6yo0n
wJdzyM7dSj44uQGvswfhF2uJYm787E4joT71j2spfF2WRG8DwDlHFeGYlNxJ8tE4
j7td7gMlJYgE83py5CmK3wS8BSQlJrtP5pCRcZeKXYxjd7Z6fraOAPJ7lV59vr8x
sSv+qHG2i4S4PJ60KRx7cPFpTj2uLvM9DeJTWM4AblXVD9hSE8y7ufzSSWpQtDgH
0Njn3cMedL0Bb/mTCSNjwUFEmfv/6pkq5v0VKMR6Ol0yHjcrTHdqFLk7ln9f9hVO
gLHkLoieBVzZCeI2nB4f9sgvGodn9H5ITtC24kfLUkhqYN52F0b9t5DFjeCVRD58
3SN+P4aeymFoNDr9t5JQyeAdMBVN/xm51A+ptBCR9eJiuhM3FCrup4ghcHSYK+ff
iaFopt3HihY0z7mGidaBEoHjEZV4WxzWgJIKCnY67NujIiCZZ5XFE4O98+H44WAc
tXwEXu8Dt+cwfERUBJGAq9vpyKq0Dq7OkYjkM2cpg9ZQnfWl3xcGs+zEsFK7vH30
8kkuIcLjDvqwhjO1ApNQcNzTrjchYq4npOskC7qDZBVJGxD5F9OYShvvuoPyP+bH
SP2PvXiUG3GeiQThGZGL7cgnItqHiduSk3iL9fTpFaqFLYhWetG/eky5oQGJo+gs
REBT/lgPa+eQH77J065Z0Ziyjz+QuYJo8tvDYoZf+YiEeasoB1UMd/qgKrN4ZYYT
zjfwKcY5WY2Ftd9SDOSw3SG1D0EuYlulRs0NYHfkKGBByhDbWb8Jj0WohOsRu6Lv
UG/R/YMqwC7n0zAfZ1qiEnAo494cnfcp2JLbK9bT3s4gEb0LI1hUIMVy3debHV1M
OkzT5Pu/YGC540LyXbKZWsxZLB9tofBMskOCB0Efi2M0lzah/r5vmX7543yiTcCp
FXDhzVhpIeCzEtV7n7zoXZrt/Vf8yxxlwwlBz8Hy2XZ6JWWUG12+vsoMGGQctJ4w
uY5Zj31Px39QCju2xNL9nzDhd+ep2bisD3Cr7J8ewqZmFu+daj89HrDyUJWpxIvp
Xh8ndpPtukjvHenpFi+EsC3QGu7Ztk+3gjvfH8kQ9NYGynhh7I60U0v+rF6xpkBr
MjyRcfOTtq1mbUk9g8I0u5Cd9xcuGaXCh0N6xfgtGqg2A6znvXdgT30/cPDvnotB
0JhEB0+JkYhNixBdvI0oyHIlXWgbJKb4KIMQkImseJQaWA3JMGzOYTjDry0mj4Ms
lknT76Jg6MzX/ofoZGVzsVwcohOL6qEs2cE3iPbbWiDevn/JwBIvhzHKMU+YUady
smrklEuRfLCmL7Dg+6G+WMgreAWptpTrmW/2KiQsIK8RYOMEvTAqbU6SwG4vGW15
4gEQE6pddacLkRCKupHjlmVFJhCnuVAjpUy9c8iO6ibjqhyTJXNYL11dEbZx1B5X
M7KYiW/LRMZdSONmhEWQ3ADGLjdPzu7Ym1FBL4gtZGinXnOC/mdbmV9SmGaoIKeo
jrvsy35tiIOWInnN7CHvRigFiWDn3BdU9P401bYZtE0zlVotwvj5OXCrv6ImGV81
swzDnmnxi530O2TLyaEYIhv7f6N4eblkJEY85SPVhtArac8Ez8gCb2Tzydtijlk5
Vl6HqgZ/xUIFkGY7P2QiIpby8scJi4teA+MMRSyHdVlxsuZnK4JTQN0E8iwQyFN7
8y3SdOwTsSx/K4x6KUDVMFcKT6SZ2354AwfOG2dEzHoUATVfk3Yb7BT5vsvvvc0R
XItWQ3ZCe2nf2KjsN8GJgUhzRkhvCroCLI12bBJtf1fXgpDMQNEVLFSj6ky7wjJf
6Atz4cUoyU9UyAhrcBu9AaGm/deuNQwxMDObyZiPe9usG3XpWb2rdQIkz6pdzZqw
9t4n6GRTf0F6yjxYx1cOnGiDum1eVJZdqpdoCx41j59eB+OZZwT1gvgoDC4GEFJs
9Uf+DnVZOfQv/1182mcHCevKeMgsn3t1NOU3uJpa3B+00kru7plf5lZzxXSTQLlD
RunLMfILo8ylTHWmuxrib6/us/TYKF3ZnABAc+RuOwY99qpFz7oP8vQs/X3/wW0U
7HRpSDTBvhSpz4NjvgbU6jC0W5l7xA5Jl7EgcKvWjBHiYb4HIaJ60DJ/1XKYRVJD
TydCfilUxt+Tq56RATXSLtZXCf615W5DitfWUmp7mMoFd3+E32l1yRlhPWXE2PeF
p2UioEuhPsz2j282D92ogoVE5UlM8cTnJabwnKl5q8v+hj0vrxttVZAPhHhvp9Tn
fZo7XYJtbSp5fK4mkx9b/l0T+1HNNqtSu3GZ7R6JibOBjH+CbbpxtSPgmA6tqlgP
5wVJhs0hVeA8rcEdrSdzuIIJ+VoQQmSGSvj+PlTjYxMXVVQD7X41eS2vN414bKw6
gWzE1wRvqKhGGtS88aMg5tQv6F3CRs9Pj7JYWWXJL7yaXsSch+zN/fciWJl/NvbG
6pk0YP4WJpaSpW4W3F1JaU//Gaoknph9xt9Y8ViJdzuaAE+sko7QM8jfQyEjVxgf
2ZcteQLH/gx+NeLgb3Wa3R/zr1EsAMfgeWl2g/J/St7GtU3MBtInoHd7UmKztI6V
soILSnHsBL2ssaGEEDc+p0c5Gb5p0ji8ExFwsy37rjqBxcwNBW7VhXAjCYhd6YcU
Ejmt54Bq1nFtamoxAop3clhUiug36MD026kMgihIIHlbQe152HGBBLhCwmM0X41U
P4i3PnOukvJEwtd7t8hE2l5MYEunNdPxddp9BcwzjTQrJHkoXTjgUSC30uhxQoCm
K6g9f5YRhSYa1iWcZvnHHso0oWoi0tF3XbWZkt/1llK1gsUkN211j04/J9PYZnfw
3mnJkFFJAMY/EkzMTIdPcfTwl7bPf1CwBVCGszbv6YbRjlbRhV5osFv9Y8863zaI
WS7e3CkimPx7LEFs+Enn/ke44Xzm9IYatHo06O+t9V8igy6IlNk+QeTpKTqqgHUm
sj4WTffo7IAxiHYZcVlRo9BIOx9bGomLUWY2fWjN/zNs4rJAzl2gR/UfcGt/itEh
hcIob3WjIRqnObNK5lLZI87ZdAk/I/KetU17EmTzHeljcwg6pPTJghP//14W0V+u
UkgQqTGYtI9QWTaK62wOZwbV/2cIRfEatvyeScvOz/VwvypNWCiu7S6Vdknb/e/z
0upa6lVPiAWibgw0fmS9/tr5bEtEVEHMq3sHCz69arcxoJ3SLrpGO18NMAz14Uv2
W1Boia95hMfIr8tcR6xS7odkw3gEEgzjQWWPHWAORwelLc6EZ6rTBX5CxRT/nnId
/ReOM7Q90LlxBOYD2ss8ElHo+TaG18ZMBWZzPg8xkARh9AIysHPZFg/wa9dsnXk1
Zolcv6YL+kQY1/UW86mD1GEllQmROm8bT22t9tvrXD94Mc+mYScpahvSv+oOTA85
gApf1Nm8ikrznVORZ4Ygg1l1ZWolYABUTYz3JMgypxdVYil9f3Yi4H9z1Nr8kGk4
wTsprUDuY42T2irjaMBYG8YXlnVURHz73sl2iHIjtsE5GFjILy4B7cSy60NVFZvp
tUUerGAPspSbrfZUpVfoe2Ibz8W4i6k+ddFB8R+wlRwVyCrfGkATexBgGyNEHFb2
wXBRtzLmiqFcXY1TWBLlI+tS28bHDcciTIhIQyoDPUMScVkk8XrvbDog+BS4/FBz
hZO0P2iiJxbsHxAoBea0cz/GR3q5iNwoL2Fo+xa2DQr81alYZ6BI6XfysLVyMkEf
EMrp/lWGkIGu7bQcwmv9nbu2OgNofRfeIvPtZNLosbAui9h+EMtJri3+Yip6lIoK
xOdW/bN0GZ1ikjBg4kKM3hF/WT6T2JR+pvOnmvOw/V1yV3luJ+p1UCQg6Wz3nt5E
swYtvoCXOVvfxs14Fa5sfH/kWYbr1iMUw60Pj5YgtBzqdMNwSFTYQEBL3jTDXarD
t90L+PEBmWr/1CX+ZwjojPSnNhTz3mhSDmwNEgoLx7fe6zO8JCu193Xf67AZkDgU
V6MP5AOBZe+GurZ5arR3e5WhsJoaWdqif3gfhR37tKWitQ81j4h9dvShZ9i3jfDH
YxzyWAn4frnaHsE5gC7vujAULdBGL9JEqQAmUbl7UjBAnwAmrkrhC4njCUrVIqct
a2WqA0/hwvJ4n+0rJoAWxWau8G9pW1OeJNhCNXWCLAVk/dBbXkWWbBoJthvgms7a
38cCC6EcnV2+B7Z/xrq1PHsN3C8s9I2XYIXsuxGRkOzPnYjHsc3mBMMm3+Vn45Bw
uDZyswjExWk2tUSdiUI690tILv4ZH+dWAl/qEtMK/7EAOBo6VfW2tarvxx9GKua7
tq0jjwIemdg0n1+PpoFr5/t7l4tgBPZ0CfzBSEuE8nCZStPItrTF5uQv3xsyk/5x
iRD2YKQ1kxRvI7qlMMbOPMGhErvllyRYdSdybFoYbnU3heJtoqNcTq6DL5uWaTM2
uMOcMEuJh0ylOHmP2D0CW/6woEjCDuoCFpe2MKcm7GNmi8roIVhhSHC7ZSI+th4o
PJdK0k4KZhf0eNRGbBRXkGqAguRqa0jQ1jQWtgFrkosBLEsFhn85Wl7vmjfpGZdd
MXkubpvpTJfbpa6n4x+eaIktklpNqgcWrL0ISyega+kFJiZRgwpWKRhsYli9xCti
dd0eI0ichPLHjost41HOyDrC7hxoA9MGdqXafSErOnGZwe35ZvkzgubRw0r3V1rt
9eZd3EljR5GC2pbCEbh3yn6X3c7ZHFheWB2nAQEgli1DkHJ1bQslU34QkmSr5ldw
KnjKKipEcvjFZ0ZDHVAlpQLx2XsT/VxOkeKGSdpiuerMJH1XbiK4mTRiqgRBBk2a
d+Ky0tnw8A43Y0nrMghCcbihgNCKIGNXlI5ZY3MQeK2uRXAm1gb1iqb1ESxIv6bD
hPC07AonIj5LQ5H60DZ0jsuK6FVIAuHFgugxaudf1ONDROh0PFHxJ+GYXEa7jHk5
y/uv4ULLNj5HCwKdqZ+5NwC1Wv3odwNvUh86yoQpAw0HjYzLN0f2GE3ifJf9IFG/
d2LiMpL5qrUIkiNGmDTmKEd/DKXUU1FsVYfyLmkZrffemx+Cb/ESjTPBRCfbmQHD
LxR0gUkNkh1VEaCD76BQ/nfQDiTFVB16tdCVHpLT/JTV7F0BdFqG+AJsDO6gVL4g
U3P1FA0gMFsP9KkeIiV7uJHT4OPdgy4r9XJlmVyVLnuBLr2Xcptg/z/jrpB2f6K1
SeZoHcShd0nm922uNiDZdYIGbG2GqrytJepFgSGZ+MGzQE/2HbzISD2fOZXiuwg3
p4UdpGwo0DKU8RVpfY1WRAVT2AzS0+u99ghyD9YpiFV/Ms7gKM0wRZnTLTC7S1Nb
JHeagHB8c9bqssSu0J43uDz2hlc9zDlvEfQ0KzKsRUWQ+xMuc8/aqvbINrXr8d8F
f6CYYLnpuLe50E4FsCkE0SJr13iHLbH0nZhBOjtKoFxUdxjmyfX5pc+WEmRE5Ox5
D/9t7732HVvkdW9FA08NLz6IAJxjf8OXXBBUoKVDe94wQwmDO9+cBdyj4t4I+KBD
chbCjlRyNwkHeqPJgvhQBgn9quKR/AnoDwOBCiPnpEHojSgbwCyXWWKulodXJZoA
NDcsYmGCdSz37MNvQ2KmOsd0mpG7h9Z8g4Uj/OTE3PcRNUwTkHvm3/5nPYFYUXOD
hOkC42c55AvnbvP4JX02x0xWTLu+tYpnmUoEE1PCdkngpipyt4YsKct+8B5Tk6Kb
3nEQNc/XROX2JxKsaXIJCkT2S9af3/mkgRAHRuoJ5LFF+wUthe9zxwfmnPksQ1No
xRHcc28upqQuUcxhXa+gefW1IaWj+USxhbl73HJYqyFbXa/91rj/jtViYAQ8hjBm
N5hVhabPBXAF8E1VoscFBfOcomLCAdjBqQRRUEkaNQBGiY4ZGZuIFndkB1Jpt2CC
h/nOmxOjIph/tVqVg1901UWgsFHAkFeiVOAwqUorFN5MReas7NccBzo+H24tDMxp
DCF6KnRulcbUG4014n3Q1N/w4D8ffTfE4LAqmmjKrrMvqSDUDU+r4JIMAI6CXQcC
xQkn907vqqS1AqopQB0epTBfVHkcHH/1Qrb4ZUDbzDWPRIG4fG0dJt6F9Lceeahk
OfSlEUyAGoTTSU5P5h5X6AavLG6AJZwr3Ri9FeDNwzAqn7cORzL6NGRaPc3OI0CX
QHWzqplEDTrrv8ob8xz6HSfqgS8p/eXtFYNjjWpJSG6mD5Z35PcjaOVcPDob4k7d
GxZRlhU6PFwM1OP8xLRwHKDZikia19gSUPD+7+HBEWwT1igB6RWhI1aVuPxHZiQA
iy+n6Cfqijv7iciep4t2GdXHfECdZ6734sqHTD43PBB0THaE7QmxTjg5l61ppBbl
a3/sd81t1O/tnFi76FrvqlyXdjZ/LqZ2gVzcPK+oBAqEHotM6E9a/pMPOcXq7RLt
+QzfDe/ml0lvX0VwI9bHffHY4ZfYsj+TCYzuCDTkEcHXYhdaUaW0mCqkaZZhWv9T
hoOetarDrFYYO5rF4pMZmfF5x8ydTzxEO8qkM26JteXXP51SCthwpeRCKrq22h7w
X5/YiLjoCfoCfPuLMqlkcUs/oqntOC0wJ/RSkfQH9UjfCf51fDcCax1bQ9oUY95S
qM8MZpAj0vb8gZyc2DMfbfsJboua9EdxBxXEVXXiw5tehfjahQ8xgtE5J4sevZNu
oy0P98tY9QmLiHV0358teJiGSq0mIwnzeysgrDfxaBmRmrNsU7ZiKlkpJSBBdUp8
eHbjUEjMCElRgCubl2XUIJ1rsjGz1Lj2Wni8DdAPqOSvPP+hVcegoXUOQkES25Wg
SzxmAlkByiKg3BcjL+38DmVMNq4+otECMjo7QvDYqvxS2dwNgk1JA76aqpJi4B01
bhexSiXZ4VnLqYPg0m0ebpV7XeIfzL01oEFQB+ya9kTbWxNKfoivy9zYrmMMNGnu
9wT74KUS30Y55m2gYOtYCKZdlwCy7YlmQK/aYFK3yAOo6fdvEr7f58q9jysmMwPX
mklOj2i0ZwsstSPzY0QnYXFpJ9vVVPX/Vbpt8a+VRdfd4FZuFY6lifJE5oKXmwf4
xjL0ndgWPVSvYlCc4VY8Amm43AXg86p7evmRLLz2fV6RtyVRvAqelYpDB30MZFo7
vlnUA3E0VpZ9BvIV6SJRAp/hUgpbaJk3i2z71vRb3bWvbHq22xhaHnheUqyo7RKh
3q5e7N5Vo4CXPa4Yg07gxFpQtlAm2TcN+G7gte4zCk3jJU0Bl42rBh/6pKgGW+pA
7oLPLY97BQSbV1sM4LnTKhsv+wo+Zxiq/DpsfFomT25x/yzBs+UbeaqhX8s8zZky
XnTSKiqV3ufOPPEFEMCpPFRFJg7NKpil37NCZxu2abwPNzU3+6D1mV0DXvHAsU6O
CUZ4qSVNCWULtLSEsCHEiSUN17u9rvF1zsubsCL4q5nFp3FzfU5PCf0iF2RhQk5E
k/ytoCLi9yc/czF3s7GHll9ghOCsWLRJllRfe/Dd77L9SkjyelVtYBXFznCTe+9x
v1dpyOXpNKkmYOj6EAYZZ8GUFidfz5QPWfpFQV6wd4ho1riLb87h1CZU8hRMwJz8
PabbqaenxDnLwvTZVtyzL04i2iMFz/KNsx5UvZImEcedLoTD3k2kGjbo4JNOtsWw
suMUJnB+E5emnBisRu7GSuRpZKluK/SvGeU49vUe+ytzxr0us8Z1EYTSlXV2c24v
RgWKeaeoFJE3B2coKVyt4ipkoxbR0eghA0PLtVurQWRtmTgGhkSnlazXOSvurQOB
FNUIelBQSxu/ERa7QF2IFbMuVWreFcT/DazkF7Pjm3oJg3GRcSZc5axA37cqD1pr
2irOBi7VMk3qtg3e0RQDzZOl08MhajvWmMhdRH+w8GkpxDjOCVKQH27xNeyQCRw6
+CxI0G3avyrka6khk9jDmAJ7fns6cLlpJQGXeT5THPe4fDnkzTCZ1pkoyAhnz6an
gp4ZZkvNFLHh6kZoDcckRrLOosGylsynccZqHMqtqUBtvtArXX2d0KKYWBNe3NA7
hTApDBTvQ2ZGtjHPwvxt16lI1k27SZXjaAHsjXcAgB6jSpfMrcUJtBzS/FrzQM2z
H1XRuPI7FjXc2YBBmqjR8DCNRjE4hNsbQzcebiCYLZZfV1dVcAI+sJMq+rs0RFCq
phYUNz3VvspmwK5quctBgYv2WUng/OzstD7zAE48n6xRhraYNC5wcW9WgO9k7YLc
g80HEr4XPQTJZy+rSc+5nVz+4EPenPobCRZQkezp9gqqg4Nayn7shBSPHvoeecIG
3zGQdK8sY41qnbJ23xiJ2YwLlHIKcyFW0WwFtRxD5swcsV00YHFBHlsdnhBT5mwn
VK5/iczLh/PjCTPZ/vssqZCEbs1l1XEnRuANaRLA1brc9nFTl6sG5IVpP40OjyYF
E7oxgd5hX74ApDAqAAvJQCgufxVBjtFr7/dwgAD0rQSLEDNXBCBgvKPkYUMgPREE
gUslCqNBxoWUorDF0MnzUmdgRKgENfmZe9eI7Z2LIzDFGviPpgNQRQhAk2AkZXEi
cDrBXlYXcOE+883kv/rztXX/7GwMKxqHnz7lxy1wN65KzwHs+3OMbpQDhxD3lLmQ
XwJBgjMKiWZYnwd0QroN/zBzb/QKCHcSvyQmq15eWoOCuZiMhCHhj1zXBiH4JWwR
tobCJTpYsvsAZ0hNF7ObIYbRdRrRbmoAC2d/FixjpCuv+fn3gGfiMPAAo96Wnc/I
9txqdYVv1RtnvobaqbDXmNVBIGne5hPExFlsLIrSoFN9gpAHXgfZ/Zi56V+FWl/i
73LSruU9wElq6BmIqHs0CG2aJxvUA5TCs5XTPaZ2ApGQmMDDUc95B2wJdA/Cl54H
h92Kbu3XAEk47IoFAjad8n4PBpHhi5nIow+V2+jEk/LbEECK9uPaNc8McDt5c2of
LNAp0xHTG+MUfIvoVxa5EtlBCQMxZcN9uw4F+0y/ig68KwmA2Xz6X+qZz7310YXl
Rx2z9aWr4RrklkkQlzKIwH2oOybhG7nWC+GjoADQSS6D3OE9nJ4T8nzZ7urmuKJZ
wX8P25ytdVsSwnY9pKDQwD39D62bBIHmLw7V0idoPQLpU2dxPQHTxkvb+GFGZz4C
iEK1crKc7j1NIfThHoo08d/an8kOQ5Tscwo1j+WOa19zdr5F4QIOOZxRBnUbq7DZ
Zu4xVOLzcX15qn1wPzphnQ/msm0+gDcAXRYbSdWQwJsFa0XnF2tu9ljcAW/nas0n
lvn0aS/T1s8R9UZY8plJjqCWCBUJkEiitDmqZxIZ6F5U267vG2W1RVh+/hNgaYM/
rFPyQL0poYJMOX4jFD42KeRZsK0eZ2pp9e52Q7E8NY6a5rcSxaO+rUrNJPjR6/I+
zAdJXljM+X3CxErF0IWQAmkMGNrDJIU+MdNwN5nR55MD8KzWEfn2Arxqgxe94Yoy
DBiu3axiF/NJ4kxpkDyACvmWUqj6zVUHWyozPl3V4Ln0e/W9wMz6x5qKiIsehoIk
4ahbDsze6op8zQYJWZTiIhpuMTm38A7+ofcenLuSLMOE+GMDUuBykZSanrhrTxd0
v791P8VyokXISMI8Z5KFBfjfOTdGV4y+QWKh2XGzhnvrxqDdPEO97zqnIGtStxwZ
EpaJwgqdL9SzCcVu9Xh82gm6GkLvUlCw7rS/Ur+F8SHbnZTp4UGHOk3aRS5Ozf0j
21jFzIWvbZWedkoSS2bcBT5YJIemWW4zRozMkzGw2vlRr3QFZYRC+wh5VReyeJwc
9J+PxCqMuwtJDik/PP9H7iJ2d3fRzLYrfT5QKCMOqIIDVHfLwKFagtus9SuFBPbR
c6alYCyc1Kcnq6TzdGPBkjHWCOKjRiLbK4pZl1X0K1RCv1NjB/8EKA4LkV0wmsle
QCzZRFOdwso5DifTM7OY5MaNAUPaUA59sg8Q5aniz7VoaMot8PgIGFRSc3GF9ynF
7QXlLYE5CRMt43iny/MRjpjwksX/Cfy8lCGU2Ok3w4oh+rJj1/IN4OfmJRCv3fPU
KsZHKqovSCg8Z2U0aQuDNH6g+J7JBhJrB9TgMrPQkW+LiFRunR2HopRSeY2NtxLK
fyuR84fYOjOSIDzFfUa8rAgCGnjLvGfs/aaaTz+sA0YM4t66kvDaF1Ikp5KrTsR2
StVbNco5rBXdzItK1YHFHnJwJIEqUzWL1xzm2dzcSBtPpVbP/m/NDHy4V7jE7C1u
vxWb+mO+sFQPzjnjZ5ZPGQodE8tGtsh+4HW9dFMaV4Dal2M/2jNzAl/9lQh2Kzqs
nam54eVqQ4UQuBkEU54cHM4CAszGzxGHfYxQhsN0t57jSS0O8xXOKVHnuJjmJj2G
jCVV5lg79LzXuVi+cJYoCyGusqAGxsZp87iW98iMv7c/Hh6TqwN47fkr7tY0ea9z
349+06LLWCEXc3jUROyxKpT5A0aFqhe6LVAF/GiFBUotY5upgH1y3Pyq4ZRbsDlt
Y84t52vqBLoCbBn4vPQGDW5NcpXV1wNSDqjdR2gdc5RZdq/qalxVQaSyl7JcGI3V
0czwUMio9YpCelLc8Ac+9pmTIOu3Sp6TXasoCf7qDW1MATIazMmUNpMgFS8ROyKp
E5EhLb7PplU6vvOewgxAF0RG5NMHnCSOSyJPV3mtEEaYEzH0vGQ5eb8kCSL2AYfq
O1PxuntEYtu7Wpey2mZGLx4gj/7HZvF0fMzWeHp1JJXaPJvNMRZUYF/IO4821oai
37rMp4FqTuqAFS/DnbBaJPvPIg59qHmh7ss27A1sr94nFKJ0Zs2Vmbt+4RmB3Cjb
jd13k/kvbZbPSdB2P+TS59S+fHCj1HPdeW7rueCG5SGMCxsF82m4yM0tgx4gqJfK
o6GtKGkksGbfmPIkn867iwOGUZYy2J51+lcMFKN3kUy78prxF6vdKDQA6dybgZP1
zfpGa6HFPY3E0bmX0HUhDJ0Y/FR64G9FJQ3HHFT9S2k2kBbEtPodDDQckfRcf4tA
UHEbnZtedju1Ylfd1t9dPlOcjO88JwCtcZwFUYsURtfu5H3Ab4Sq52IZF8GoBrdR
mExKGOCbvFLTWZox4gL0eOjIvjJv1Bu4wx//H/zFzd1jYv9oK+xlbL6p1qZuJbD3
uFWleCSh+XoZPKVFFR7nhXkOhI1HF+8RVFIha2aYazYBGjmpN/xBzGcccZ7S6W86
Nfxp8o2eaOrAbm+7pqBAxuFxcMlbTMRIDHxREU2uCehju4m1pz4mauoRSg9GRjPc
BtxR182AfSTeLJyIwf6k8l2sngElipgqJbfDsu4UvYqKstzJ9gDWPOufxHphlFk6
3EjnulybyBCr8TCAsI1JGt3rCOIek71Hr2HHBNSfrv809uDHxia9JT3GYEp5gGjx
GInVYdK7eq//VTTHviPiODzJpEQp5Jjhd1UPM8i28dSodCoITXF1g3HQUxXkuC5b
rJ5TiOwRHsXZdUUBlukQS2/KXOyVzBmExpsw4PufI+BqaWcxoEb06aGuZIDVEhKt
uQkhzvpFT0ig9DdwD7Bee6P5TljogGanA2GdbgCvKeBA27jY7Z/21Mb/a+RUYR4v
bJ1xGLEbmvqyzI6GllqY0p3btls9E7nEpP92wjX8EJK2sqO87C8pan5qPDtLS/Kg
i6guSRnJUOvuJubzDvhFkUAqHkd9Q33jhhGOHTFAFHLaxmLM/VfxuG+PCzUcCMAs
zc7dOWEV1TQ5HtaPC2Gn/VQPHOC5wP1TPV5xfsZ8rqVWgiAbv+IiJcUiVo7z8hGc
5hWQdaZud5fetWbYQ3O07v3yhAnRDJpN1CwNsEBjLDQ8tt9VGoT2CgWSVkssdZDT
CoHMuVnYsbWTIVcKhKspz7qISofYt4yXYBEiq5yjMHmoJ408jj4rkb5rQ2ssu7o9
ESn40fa6ne9vBwn2TQ1yR8+U0CH1EQ9ywHF9xyqSc7bgruBTwEGe0cYQqAi+Ix1K
SECkdWkSbYmWYexqS25Oy3qnL0Q7NS0LP+cs7x0rXyhzSvUHJHWA6OUPlPbjhmOK
MK4pYTGpG5D1mAUOY8t2dt9o7zinK2uUirmAGwiJzB8g0/zWiLp4JixMpZaJNJlA
l5OPzUdt23E0BLiEQIn7zWdyOpmPM3GksJysMKt8HOyi3CPtSCOCKoqw+9xsWLSS
pu9v9PeyXOuCTRwQitlqMCXXWK8r4OAbguLtBWsvMyn3nGBSV1WVdP0ZFh1LAy0Q
GXECjrNoehEgMIMDmh0vKayqJEwwxCeNEnLaq823suJswV3UC8WJ1lK6+1uPgyP6
rKhkaj3w8D+WExZh95mSnZ2D7tVZ8kbrYEZ9gL6FKS26D/VN36OIp4MsWh1XOjCT
xkUuZvmd9Nhnv0AKtJldAtD4Pgo9zCjzdoJKhxRJbI1fi2F3n213LLKBn5KYxXoX
cN2RmlLe7edIlEayh3Kg/OXM3laTIC31Krj6vWdrU5srOOq5s8KM2MI5E3xCPgtK
zQGNODS3HuvYNKAsC3NtY+YyZF4EQRTZ2Gr0eXl7PrvGm4uqCKt1m0D77wUNiXxa
AKNT+Zt4PXSbYiSrRY7L64fHdcKHmowRzOLUILERvKlQuf1JSg4FIbbAzZPcTQQw
cFvM0AukllQoFWagu/KgNT2Yex4KAgODIsQxVWxect9pe1axT70s62qzTa9LAEp6
ODBkTSWz3UlBeOacUrcrhj31ytc3wQTGHMgEkpcYtboA8IBpIZbEr6eaYA/sn+WQ
q1vermHm8pDgnHrsTeuLYiKWtqFTDvne6jItt8nIkm896vBlJ9IxbLmBOaoFC2pb
ZoCN0ZKWjGa1tclzz0Qhw9hrr0cRoizMaKFIFmtHS0nKdqM6qXvsA6wlogAD3beh
e/ZpXoWmvEzcOO7rG7ThYB5wkTf3tU/dUwkWMhMIJkDgO8rfMIS2tdRhxUQ2JS1H
NoQHDvhjbefJ1x6uEQ9c1u4BMPHhBrZlyw1duxw8PoDuVKL8GZlZWnyqjH2llnFX
9enzb/zggK9GYVeWKmd7ZhDrnvmgT4szhj117RZCVo4CxFy0xk4fNSLFcLPOVxxT
ewUHsOsajPwMEVRkCoRF1gZboUBTEnDhX8gaVpOgnceMXtaDkqOhc5TRceeNF6IX
qw6DYuiA0FAD5GdSN5ANT2Vx8nMxvJWRkkoil0V2ia9dTSMj2pMphZ7Zw95lKW0Q
9BmGysCeLaG9vjNszNLxsVQ2oo7NVHP68a7kG5iSjS7jTdNAUOVx+Edr4Fd7YhEH
4RBUcHX4bppiQUet8430H24KM2nz0vkXi6hxi/LVJOvJMXgB/42JLwbSYXuBLgFV
I6A3qaV2cAy/llaEhja2TOHXIjwrH4cADQSRX1CiBpCv5TzU+2VzGDu/97ZsWAqH
SMPZQoA8ztkn+pJmcEiYCCxIG+I7gwiN1eIO/0gY90wOUnU02xU8xpJKs88zYVBg
SedONSlU/iUqe9mvdpX+ibrmkZ6FxXl9jUN/COkoLHJTBWC4ZISNeA4NsLNKdWTQ
Sx9maJGF10oJ7VMcA4lP4QeUOtR/ioFAndTxhZdeG63Rw6cWuWgX8a+zslVAVOnK
TK8gtrgYpQ/9QGvTaSfooPaDuQ5YgRgVBgPbJO2m+1ALeFKHLmwy9qQ+SyL474zI
BmN08z/8C57Z854c6DcJGUCmttVwUF9lBHqZJY6IFmllx8cvpkaoWLdFvcTb86ff
i+MKkDlZAhu1kdJa8ZsAbjJaV7kR/Dv6XYJ9w43+idROB4uWhojv7rUVCbVk+Mr6
29KRTN9BErbDIal1KtgLIjhK9m2p6FoEIsj0GvlyjfJZ4FxgAy4zlfwcAfhTP3C7
r3ql6DUyIAOVo1ELkhm5HTwLcXtEUSbenNdAq+ew3ill4TMbzhB2Epwc5vONAn74
JECD+E7HhOK8XsQXK6ZyQasUdRudLGv00TmcPx96xduHYNDTkjwX9bohtsfdX+9z
1X574tdwYYBEa4hcfraGcD+eTuHC3LwxcbEG+WrFZiNlwRwo2fnJxwXOXdqDDphq
gidqQ9++ViAEoHomKWKTIX1DBC8ugP9gSehvO3aBTWUTdhlYgg7wHG5qeFBZfae3
WlmpHe7fiYPUlm9DOQZiPYjaKLHvqISKgE0Cl/hqkpm/GzW0qNjvTW/7aiQhnYpV
YYFYosq4jXiL/fO4lJP+cePdmiTBabuOQHjE7h4RG8khVVEeTJzBNuO0yprGkPvb
PbIQRZAKDV88Yzx1thaA+JLIk28okaZg8qbMsQ/XyIhSVttUXAbJjzNKyVCONSYR
WPDCfHxTonJIn+WiHpmFcycDXV1Ebda/9tr64qid370pUtff6t76Dm+PNxHo+VZ1
G4HQ4InnTVQ/+3amxibRtaPeyjpb8EvWKvOLRgMwRca/wWiX6FyGYhzIPcAIoeBS
VdA4y1iS74NPoua5XXNuxO+aC40Ewh+KCA5iDDN/mQfrhVd2iFEJmXNxmtQuctHF
s23IxOKDzJuUgP5myRpm3rciZODM9f3wIzwrCEVGap9Y732cyY14ueCjOtKqvABf
JdhjvU681SvLhxC+QTwIW5CTzHFeL0F9gcbgTELjs8xWLn+H4gE77W9PhesJmyp3
2gHOZbPCTBQ7uarfp+3XvBcfLQBJuHwNkDs3UyY7o9d91UgVRlY2QPKtASjxFdPd
xgQHW+yUX2twQq0j6jYc1/oUkYA1jnHu4HuWYGCfo0Y9Dzh0jDGy2D6UE/EsKoE1
zkcWVyQSzOIx8GML1lUCkJ4aOef/Jx26KOZqXFZBA1DCLteV02MuExnbkfv0luwk
BhfDcocwJjageh6anio61dAtSFDXqfGFg7p8PM4tk5Eph08UWT8NWSUF0NsXanCA
9G7O8WQriFYeNNfmjvm16jELRm5cdPIffUecxd1JpgUaQWgzEzgHiIGrqgnJFeHk
svH+1qb8eV8v/x5c/2qj2L8MwEjZy6fd9aEbOw1L8ou5KjslnV2jaJsFWcMarcqq
8qDUhbcrErPizPe4+v69tcTLXmmbJHuOeUXVZz7L201B2jEFMFADqNO5U/ShUNub
zjxfzzdtDm1zi58cba+LW0egRau5H1bQPhK6SZiTuwel8WCguR2qG48z6KACJxxd
N3kNc/KCprr45jMd4Nt+hI3J4lqamUKK32clsIjH98yimDwSeU85NdjEm2BT0hr4
2FzC8DD3V46NtRGmd55cskyCQQoXkcvsmhbBdsNgMaPfGgAjZqCoqaZHX3C5wqvo
y7fAthAaY3GtDti/2SVbt1cfwThEgjdRQ1c/goxIe3KDgNOzEfNrZwLRpecE3+Bi
cp0NE6GAiupcFgvFMiDAWSKbLZNVssTM6qFP6vW0rCLj9HS1feyLMh5MkDD8OYa3
0dLZea1W9w3UUKO2T7rD/2cGChgBWg7Cu9ZHWqNZMHTSTMeIKPPWKMdjBU24/fIQ
9Jwh0y7dTlLY4jpYbbXl7bAcETaVuie4uVchC9xTTS0KeuQ/dxXEe6cZwSY5Uf44
kSVbAZi6mmaNglVulwIFonr26Nwbok9t2VH2OzjQk8QDrwJHANbCojVkGuUO+wOx
M9L9BFdgjwxxKAiB3jr2scM1nDI7swhHi9+NmLH1M2R7nfKZ8HnwxK6De4NzhyYL
W308zwkLDJIYnMojXz0d7P7bUfVFvybnSZ7h+o4Wni88u7L65HFO3ItnmmCIwP6j
KQz8iIPvEEdGJV1cqNpXiz1/YrtNVT6IbHpgfXlDaefOtktVy6NuQQjHHKjrXSVt
zmYHqoX7CtnesRP3wnx79bNFde95h8ioL1lxjAb/JYcDreL4OqmksvHhGb77IET5
SxpOHaHar2khrR/QOyyHFPieu5X+p0Dd+ZjHDLTDFW6yuufMYJKSm7qGzj8qypBx
EetS6XDN9QmS1EwcV9LjZpj/d9vWcEsAWEd2Lpf6UCtRcKg4m+NQ72mizVGGDZgq
GvYolOKNCTSUSTa4Y6VUEGfcAtT7Ol2ElAVtcu+vj8PtYOhVyFmv+lFiVlgQBKUg
VPGMHHYhIXuiuR9dchJjyTmilBvi0sIgLRnKHN1vbABXbHlhwcyVMkUDNHNyc0V6
sQqJHMtxAZQIxeOO58miGO72RzSJwcSnOuhWt6HnpyJoYalMmhhW6SLcnHsqsl5Z
nLfwmepfPr356qNFhW3S1Ix2qAkJ6opVUlaR5sqajS/O+Y7M067GP9nKSZr01FAO
/GP1c9uipgSWjG6QZ5/yo46nSi1qC8Z/qByD+fAmwPt1sBm8CsoDX/VrnjbOVQ6l
Evpse6pb/eDLSyLcajxeqTObpRCd5s3dVGg0OH4QCgH833LOjGWnI6VGVjdv4Q6m
gJGiACmOm+DKeNyiBSCXAFykdO+Lv8VO54C0rJeECLoS6yIW+mqgQHW4QKjnbbCW
2sFMi0aV2XGX7xjGaCzL+AB7h0KWf/yoW5LIOMDs11ohPF4exVUCg688iHT7QTpz
G9r9YYTNWnZttj2gJPHkKOMzvXF8e6Xmy16ethNGrDXc7NIaBv+/44h5sHRn15zm
Wh54cUElAvI6rFh2MlwOceFV0NX1lxsT3jkJzAAw4Skr+h0ixThoaqTOTdDBXoEN
6HHauGkFs6qpWKmA2+pnnYwGaWEmkuq1bNFrnwlqyvGd1acVIJvtQgXVj/CUxspj
C+gLcFpxxkghp4OlDB37jM08qoIfGOdWBdGIyTAEXDGTyarUGDJUbhuF4UxFN4x4
yyWukbA3V4j8+e0HH4gpWcyVDoBnZMVHoHlziYMdsvp+SLtttnmxmmFC6GOJdylB
fyiurpncUGFemv+MtwIGO1EEgXYlvGF4oIOinrRMiUqwE4r9fyB8T8qJNZyNUWDl
n1kxA3K1WO0reOpLwo3U4IibPQKMxI44Uzy+56Yf8aypxhOh9NUyOO52MEG76MwW
SuvvOossSkEgYskDTMIdzkq9hxJUfZDJM0+k5NzW8cC5rHVe7gcAzhhxvrZV14XZ
cs+kHwnyKJSHy3RPoRPptoUtHr80/JSr7ZxPukCpKLTTSlC+zygVcKAQlkPFPmPo
+I3lpC0MC3r2lP4hrxkb0m4GUr5QpctzmfT6GOZDwrqtRDaorN7AX5gXG3c8/pxe
LFefRaiUaALEJuVm+mexl3i8ndoyXj1/a8zxCOGHtvpCGp8zEhslIuokyLeofxJ3
yDKkUzjSTFc+9x9tBrcOPnjjzB5nRcbfmHAjMQbD+AIepUycV8xmgFFxqp5YQiVD
6l29PNvv9LE5L1Yrx3bZf9c3DbYj2VTthCJRXpX9Zblo5D/CRLyF/pGcwn0FBDPA
zgUzQOwc8K0rs3TE0zE+ZSivyEKHOI+/JFGuo7wbB2uv26Xbl1Okc/JaGXM02DoX
j7UtQPgQdgYoJv+PYr49kB6ZK8EscaOZBzP5Nzvh26j1Kbfh2m3wJfwQR8fb10Og
eGmvyM2Tsi17tO9xcEmWBf17IT2d3QwNJ+pxfHAKoI6VIguS40Wiz0Cd4usX+uIn
56a77jquIq/M+pKyyvHDZ/6XNm8lRypfkwNYrue5mSk3tKTOgESl46Z0O+cqFBNq
hTb7HY3Hd9LqdLVF1gmgDBmIXf+7ctqpfBbTMBXLigyAygWjsXUxMeePc/stv/6t
7uIu9RI1FZxW8XfswUxHdBEgxz+n81kZChzLrHxSrMxi2rZba/jO6j7jR4Fp14A/
oJsCVJkmILjkvGbNho28ljJ1GV8WDR3vmnZtmlQNiZcDEoa4YNMiNMtgUn9R/eaH
Ge6ClZTVTemTbQvKWdfhf8BWaBvzTwwzyjlBrzJZOLA/pncTJmrbpvw3HxO87e8s
9IqmMJO75JAKfxb5fRIWlYNTDvORWt2BDuDXUtGC97ZFR8LVD0+OzuPWDBUIyoIS
AavHBOq5oOE6B3ykeqsnVHeqz6kNWgYvTUa4H5yuYgOLwpR3rFvmoRy4axLG5/oI
vH7zz0rAMVVowGsFVNzO3Pfham+GkRZ3Yqou7sA0F7Ibk1VudI8OKwomJgdv7Nlv
8M8o44OqAoBiAxJhEpp2KIF9Fe3dYN0Svd7cUYwWkq8Z3ZT0Yih/L2gxMmUJXDxz
qbFUY+p2AX+Jlc+Q7VchEl7Z0/tFmRZSKHP6wAx1n05zqvT/1YR7FkoPKUKTwkQP
gj0ai9vg0Yz9cf/GgoG2GzOHHBtd0S+pyXsfZudDUGJRGQ7FLPBeDjwcYhnm67EE
cZ0p34Kwdn8L0o0LN4S+K2z3zpKr/S5aNNP9z1wu4ZN2/eu3neYQc1r7rLtonnDT
LGEBWzqE0p2d5K/SwrIIqTFIoyJIicN3tymxUoL2Oy6VFjD4rSY5qWBmn1hTONDv
svHDrZL6zE9JkYaQxSTLWzxP6Jl1ahFEuOKhctv7Mk15NGPz3ljlo8PFjNoAXqWK
SXlL3WGSjx7UnmVmLGg/1Z3gtRbGD9PJAzrV+/8S5CMYVqTbYxM0+Kw9NJbE9bdC
cjR1P1NL5Z55DfDsTVCyl6A6Q+cLIeQ06vh4nX5Oq1GK3HA5XzaAjim6L0Ah/Yjl
gjqDSsYOLqtGUWYNqT6+HajULNw3MEJt24Pa6sGid3BadR8r+MJ/diGbv/aqZ8mK
LloJjSYp9FIUFj/iOqyyymExHo8bvCn3CL12UbKjSsVZpNwPU7QMGbRLVxHj+XM8

//pragma protect end_data_block
//pragma protect digest_block
WI4TFGLMnr0CeCTfcP2vYhg9iSA=
//pragma protect end_digest_block
//pragma protect end_protected
