//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
BywACjJZpQnklF6ttLt+NNO+QY94tjxTYKbHLffzO41f1laOZ5x0Cx1kyvNj1Nqh
FtozV2zgIuwRhIxQs11HJocC2XGLV9G6oUa2lXYkLsP2REfdlpp/IkN6LKduH12s
/EcKYO/GA6pd0IuFoXguP15W/D5CbPonDP1Z9vzaiGN56hWpTRDSKA==
//pragma protect end_key_block
//pragma protect digest_block
XKECqZ2BgKh0uB8FJF4FH0HYaVk=
//pragma protect end_digest_block
//pragma protect data_block
cP4aLr4Htnk94nVKD/2NlGpGEOSUWtkzd/ueUwIEClsDumjmoiA8IsIjwObHDC8a
PRbn2nQXN54E/IicQzWOonGNy4BYWNj4qPJG6Bp+VXk5E+HHPqvA5iepPAHYoxLG
PSnCVGgAatB2XAGT9bTVYBqFdf4KQ90DaJT0CJZn+P3BKO8ELro9KZ1RP7RYMd1T
kTxHv/c5xbW9xoR5DtdpEr8qG9AWVFYCrkiCS164E9sCCSmpvdxqqIiOpBvfL8ka
1kjm6J+N3re77w6M8erXpFMYOfsnk4zhiB2pz9foNOxAtPP5DD0LsRvGaGnlWJl4
HFVvz2A0u2T7f4t/oQ8eww==
//pragma protect end_data_block
//pragma protect digest_block
+Sqg7A8OmFi5s7u3FvNHtxsSw8I=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
XBZAWYkpPx+Jtfvfn/45H5J8OuxaSD0g9wtDmx4eHUdCswfPatx5l0DyDCD5aonN
gUO9gTParFzH2R+SC49wpP5UIBSycFsgVvoKGJFXKTQGo/Tca8YUNO/xt/hRxCE1
2gVrd6hck0BpqL3T77yl25QmSWR9suSHIZn0YWW3NhKhcqQYyK0Ilw==
//pragma protect end_key_block
//pragma protect digest_block
4v45F11Csd8ZMKhs+/qspu1PPns=
//pragma protect end_digest_block
//pragma protect data_block
2zcfMOS6jZoO1OmDDgw6IS/R/ooTo4TIbRyF+D6gOwE1Q4cQuqagmJKkKlUYJh/f
eMscuYqRS6MGHIRMfWcV+rE/GAv0BdAmPvvk/BoN/70hGluVwBc4sryGSxfSAxs8
hwZEie/iFkcy75m7N6UUyFuR0UXGi0zMEAz/R/17bx3Xwhtpu+XF4el7gL3YG6jX
7AM4ZNxkLKViQAbO5Tc1aGJyhNR5JjIilyWn/XvNj7DAj9M7scDKN0/X5e04usuI
2VCbEW0QtLwU/no/remU8UfYGStBHdkvO12K8rACXdEe78ogBxAFVgGjAv9O1sBk
/zBmXt6xrle/a1HSNH8bqw==
//pragma protect end_data_block
//pragma protect digest_block
0CIV3gP5wwPIaqNrXTCht+ECtyM=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2AVirEp5JG8n622WSx+Br78+KKvTLHqPmc9gCXmhbdAqYvw9vK9YuDELM2r0G/al
JV/zxRtJVw13471MGfBjGg1reRtqqhgHXfWwsgmlgS3Xey9gwTsq3kMSdrCb992P
CRcvBbbAHnnSXHxvbO7GBXkbXFEDmlPCRo4B34UUAwFGyxAPeR6Hyg==
//pragma protect end_key_block
//pragma protect digest_block
i1kM1FrDvKfmzwTwcBqCSPtvTs8=
//pragma protect end_digest_block
//pragma protect data_block
oYXZ1ViWuwDqsaJJkoUMtIa1vLXqsNzwpqPzWrmkb02NBQrkAC1Yp/rSsubBKfwy
vYTbJwJnigbDssVA2T8/QN/IcAW88ihuE7HZt5k9pU4+TlsTVnmOZcOyzdks9yot
O70pYep3EhuKmW7N6EEf6hs6NhXSatL4xBJG41RMUeXaAwjra64tcE2JZ5SzO6wo
OG/kgt3k9eFpnjvHiAZeV/I8TDpm0JMBFRWbvzp+lDVh26b831Wuvygt3mJCu4+F
jjk+/YZ3/mnfeiUzrWZ7D6e7jzOA+FR3sZ2uJu2kuOfmwx5ZgWfa93Sx4SDTF4KP
s9b37I0n33cOaEFaYwsVSer5CYvhAllZ1ovycK24wm+QlJzVzPyU/PLDNnLYSPwc
30R8om2aQKVWmNjYcgJZdyBQ/Ll8AknVOzFutvI6bKbMSBtUfM1qNa2svIWZsnK5
frNHXxF2swF3CmoGG0S2u1ZinlIWjnuEmTyjRy312QyjBBn/9gbCfVXiyIE/Lv/3
j6RE9hSK7uvkre/jZ6hr+60jtN/w0Rwcti6FullYwYI6Rirs3haXVPh9fEVgdu3o
orgpQ1Bmmv13RUQ8aFenApddq+kdoVUL8xn45PqAMVd9ri6gA95oKBRugAqA1+T1
2SEzh7m5v4Ug+gZDSqmQKm+1yte+oBARr175kO30HKdTSa5igp4aIuW9hmtZfyjD
yoRAeQOWuSkDVO8m5TYmdBIFI5TKEZuzT//o4FQ7yKFKuFy5kkL7fKR4g60+pSC0
3DhddaVYXf5i0e6CUI+rl1gD4v/xqd5NkfY9YikIpl98KYgQh/Tp++Ir8mgyniZp
bD9cu0J7hEbkuhzcP2CRiCKMaY1KtDr8H4czxBzrZh3smV9MgVKmlYJwdB6BARkt
8tfeYhWDTRtXYFrbj4xJnMT7Ml3NVzd1evQIC0YeCjMKqqHCvq2mTHFrPatgTE0w
bn+aWOC5HYspDJkCTa+R14ZAfYi22dqxvEh3QIWLYXDrdw8/6CRBwAWz81kHElTq
++bLlVp1iIzImBEtToUDQg8LgX+x0Ypi1bGzirIiY9hyDdlQ+SIZ1ssIxNZ7aQs7
iLg8i0Cbwjs7fOrHtOiBzA4IiBvF51XBfkHdYhjHxdyE5wdW0ValFg3oVRxrhsuu
cioQfJ7sdCkcRlrCfv4wZlpY8rKsa8yCmBiT3WqCqjepjxp0jcwObR+kCDcFwjhK
Mt167EA1a5sKt6Cf7zG06UEAaaewlW8vF2GQ8JkUp9l3Tx05DmYkWEvFTjqSMSip
cWY6zTW78puFeM+0oCbVqYQh2uoYGuYoK0vnhrxse+VK9n5ERf9FbdNYRqPj7YyX
RV0FkBGYc7bba+5s7BBgbsDTLAwncAz0mhi22e8YCop0Qj3brAlTeIq8sR7kHbB7
jPNyWDlGKQioI47RnCGPu5am9OFdZKKDtHbAVPD64LqJS+ii0Vd9wttOgM7x5NTk
ydfw8hafnv37I1NVQDBRjMK8KCunJrH+OsiGb8WwtxsUrOqZxraGgr4hTs+eyePR
Uy0h1RcUu8ACgWPvysx6PFSJhO621V21RSnAZBkzUIBfJecJ7bCVu2WjNznauy6x
Wi6JsPKWLmC6DIZ1SjiGyLZfiGH4encgaip2szVJmLaNMCXjwbbhkKd97AgxpUAi
nFJzDdZ9w2fWc6/06bNLCU8o8hq1EGeg7N9b+1a5qHmKBcGaRBhLNQWDhZSO+exD
jAgOCZA/BSzURvahb8e5fAi4FknJaKpfRNhXmE+Cda4+x43EjFvCW4FkB5/bK8bh
8pgCUgbZF2VGEycD8UaYc3dgDRsqQMGKktK9OzXOednWk7vdv4cz0PeD6oggn6J8
sR9gl4sg7Z92Ac4IQzYwbhflf+jBy3omcF2P6TsxOV0GBGunNdH1yvmOIk+qJLI9
5PAvNLJarCVZ0jYk3Ujmv/7XOMnfcPWRG77y5IYanA1e7GnMWNuVogulFcg3N0WS
WwixpDaopiTHW0etBeyhMJmAumwnn/UTyuATuR4mQIp38wK9+X5shEa8HRy3T6kI
0qy2/drVBmvOUi7WLfg2Yp4qmxWpwjQz/MZ/+dOtEhPSdvVvXc6fAGs8VukxiqzJ
yJHTKzlHiRu3yV6NhRa0/rDvlEWH4kbym1TYALVxdMWeChDSXDq9QskLHj760MCS
YTEpK1ClMXPwt82e5s6d0EOlXDQyNGe+gBtoEem0bPAayYeY9RgKfqZ0KGXyUFFy
EgOUkLrpG38X3pK3tWQeMdnQaF+g8+t/Fr16M1Kv9JB+cnfWFpQv0mqjfP/J3P8o
jpXO/w/OEj9nGOWdpdQX6rhQbnLgGGZplzuFWwlKonc9GGaP7Gx8NtDrFe4jEM9b
OTaEnD9RPMK7mhS07rhuucKDlYmwlv+AJ5t16E+T00heQUeHrF//gwawR+HIjKn6
ihOjw1eeYHwCZCYV7/oUMbUjsmQNTtm+C4IcsCVC0rhm1XN57rEBj5mz6/KbzcrQ
OgdVWz6m7/byYbTMTs1jxhSjHVsYXjMfvoAomMqENAkAYUzt4vGPGvaJD6Pl7jrZ
4YpJQ62BArgwu7isObOcMjxxXpLg/j9Ts79XDLDO6rZ0C8/iqSPg3rqRR+A3M9Bp
boiY0y8dlDDAUTq54LKJUylers4tvYF/rAX6CMggoY0tkqoa+19zYMG2fSqlX87K
QhhHPTqGl8nFEhjAT3xzEUKNvdX2Hrg21vnI5zEnAGidhS40iTKTl/QP+PJUSRDy
88+Uvv2ZduIUdldnPOQ3qFlG+R23WqZ9lvmf4mfBjAcq9zXva3nzIZdIvzeiZbQl
u2y7nwuKv2xKhbCs0o8unwei/Wq3zdULYiXqxw2gcaNQhXDg6/ZI2MC8xXNiIRcy
n/XTgkdVYQwPQ8N2rwyB6C4Zl4Zk0UW/2h2FZndKK4CI4qBStSdoxr4IjgaJ0KgV
Uf5iBjWHNsytFzzeiGZvx0pdYJpNcXV/99x1kaiZWWdjCBGi2INJtrpB6Q6tgYlu
DVNT0PKI+EYVYMpiFkBJYAoNBQJT4c8Q93ebVig//rs8cTHUF5kssgG/8imveyIK
MlUCzfb2wC3G21631UNo9RmTsWYFvnTEjMYrlzEnyxD0BkQrzhTT8KoneLgOQra4
/gSEKtnC7npNKOGBeqbLfP3XIwtP6n6xCHEA5x0BoDqJrTfYhf45BnnuJY6cXcQK
XjbTOYrXp/Nlh5KKsQZ4WADgj84xxLM0HpPlvHZjnwfgkbWKPJOryucsTKznAoTE
bXsl9q2vzekOQZkl//Ie8Vk+rH7LlOlrI7k5FOLQpxfBDKgVb9p7C9o1tAS44J5t
e0blV3nGZYBDYzofjm1JfGtYkcqvoVh/By6mGm/L5z1CLY5XtuWJIbSW41LZxDX7
ZP9F90MeUO7iCcQkn6504BaOlMopu2ggUfCH8u9jMXGl8pD1fSY2z/TMd/hLtbV1
380XztcZaO1Ol4PGmAM3x6WZF6Dfl5ICNCP1JUAFOOaa8puPHGoIMk/ZmVMCVtl4
tP9ZDP6VauPWC2AfH/kFa47osDVvI/IZKwFXBz0XHzF9HT1hv+aLIevkkcaYg9yn
avAWQ1pDiqbJSAHAPcaoqlr1KedbZik6lyhCv+NN7uswBYQR+mgDQAAbzfDpGq0E
BI3bzW/JXbxAwtgeu6IRMKhmxCN911oTN8A9gB2bqhqOXSu8iQkfGxEzx+NF6pHX
IYkMIXiiJtJ6sfb3gE5ehfnXNi+PaIdaMZ51216CNLNzDeuFdQr3SSfxukk+BM0G
rCocHExaLKjpmrAQmTmTiHZ8Bfpc2r5FzMPtrdeoIunfIVaDTFX/dwVul3GyWEWt
vFM9QORBm3XP1DGspuhx7T6Hkhjqff3LVwXq7AYHlkJqSDA8oUS3BFJG6TMxs35a
xaqV0g/+dTs2H1gKGFWWbm0ee66OGXmHf5xMaG+Nxkxpk8ya/x10O0obLY6kgsyA
ez2W0ZweJ8qAyLd7B3np8BmqLXKko+ysr7eoI+IdCfZu/zgAGsqM1VQB2v4DLEPi
GO7dcsENKgHrNSV9Fb6Sw7AaX/Qt88WAhuYuS5H/7gpcociCgyo44OZV2LoU9J5A
ouPfOF0rabrRjHDsbQfLqktUWZy9B+nTn7+3+SJLJWA+FyLYxmdAO4nkRA+GZNlM
i9TnOvx/k2ntzVZ+DxiJ3dO8aulNne/kLfG7vCX+mt/+WBpt2meTgcihqsiXt802
4BNo7qBYvAvfE0FyzQg93v5TwxlhXN7VxiDJLDgAIXw+ABrQNygUdryJgiup0nIV
b87LnO6ItAdcYepjnWQHquJzrxCqjBG6aJulv/8tpBMOjC/xZPfVczwhFv7sMrhQ
EEaS+2MTaCl4GJZQ1x36iBeTYQO2WPUJX8miL20GBr74ZSOlkI7FtrNUCjMNRpR/
mqDqpho55KXwm8eVFkSn+cjWu5LBthc4I7V8Y3d61Bzu9eu3eI7oEYsPDRm5D5+W
9xkU3FNyENgsY+H7nKrf6vmImHDP8K3NkSNmXeTXgLgqU1q5DzjWLvgp67ongYGJ
+oM7C06oI11F/cLXLmRNcsWMA24p2pb61Hfj93j2HIZZQYZL4VLZezs8UTLKz17v
klCuFxbtSk87Ahh01+1E29PEy7OAoNI9gRCndhVhDv9SCzgRgm5znQhitRKNghOn
MpRISa3mXTnsUTKYs1rqtZwmuzpSSKmwVV2f4y/pDgOt1oLcGMU6q9Q5ihjZroWu
WAv4yE67nwi7NJK+tl1PmlO/OjAnqTQTCzrhraCuWcpQCW4rFVE3OhIETCWLTQqg
EerCZsBe4dGCl4j3LFE+JdakHfsRU7Ck97Eb/xgHkDt5c8jlNQWsUhHsPv1BUnIC
i5ytuV6tJsBnwBO4TWR4p2007+WdW6aOpS8eZRliQ+7YrP299MpECGNUEzWXmoEj
NGMhf+tRqRsdQu3tY+v/qo8tTwYzN0IZ5tqhWg7nNWYGIN/eeu00Dtw60eefbrB6
LIi4qKpVSEKeDof11w0jFiBfG8+/oBhvAX0lBrA6vaKhkaOzksLwOEkMSzUpm6YU
jtYAGqCxbpLrNEX4zKIfw9jPZcoh8gdd7BAAX5SeIVvz/WpZeKc9MPhsIFokTK0p
23gAG4XnsWqwx/L3fl6LTKmqmX5DnQobAIlR6+73i7m4h55pz2UsN+RGr+ILgD1U
iPRmiq1Wnq8qnA9+e9iWNUIK7fbFMaK3nM7Dpd5W2DaaT7XDhj1HViSXn2fpiBe5
BDdlmTrGgTNcXX7K+BgpVYD/eT9tlMZgam8Ok5iygsBxw4J2wNPQuq2+Hv5MvAOC
C8/lWikKPWEvmMrMVSYqwUmPT/0TWtcBYR9iaxhd5WwvGLs9IpjuTTmjGaiUTNM9
LmTY1QitqMuKLqgsM0mA4CjAcm/xyybIDgyVmaXgX5sWuvmRifhte11UPNahcdnm
Fq6ICDiAHkXZ2ydcxX2JzljAAD6jWhF8f5XMiedcCy43apAJM61iJ1bPPt+vIpg/
UqtBhvSSVR4EIQmJ87x0C1sGWsDpD3R8nptU++hZYSDITVWx/rEyUtYm1/q1leBK
fbxKJAZ+PQpYm5EeLgFYjYObdASzlCaF4W0+OclWflpYIu8bv0rp2NHnO+OS7GA2
MeTW4cHsVoVBteWaOnALjDD0xfuwj0ChNvnqG7+un8e4H6P1UAtGdsBS2tnRbVpm
ZwVJkxA1rOSJl5lCsJ86N7kS0XODptbbOfUncai/Wx4VE/W+OWPkZnfGEo0WLoJ3
5Hl45cTnWZHECSRZC3PFO09l2W3uNiHrvln9bRE52BZMfSe3iTSESfruM88IT7Ok
Asa1uUz2nz8AUAC6kcg8IbI0EdUh0b/5AWnDLmx31rLbi82MTCI/5smdyd9KI4Ty
kQkWaIU8Qq0wCFUqXwlHQa2q+0jjorxwgpEli7pWtcS/kVHckc7LEOMSBN8zorY1
6DKTCQonGvuiZfAZjxMchbr27VgGQS2fuT5gvOl0QB9jjm10YHv0wYYSPc8PZTl9
DV5t5NkzoBPU7StGykChay1jisx/a28XgIihM77urDVR3RrjryXPfwEEa9jKYMUw
tkHEPg4qMK/v2mzue7CoB1zxb1nZZUQjVej52hLLA+hwlACD0eTjfVV8b5lIGGCC
wIg4MosB1Htg7oldxshH5jjck/wvLOODr+ti2646GourI7gcEGwOX2BWus6IdV5I
0QDbpAZUX5Du3tcV7T4z9SVeONvVn/j9ipjBdlkRYmJwlB9/4875JVHLG7CQqYX1
BugYzk2GiF48kHgYmRITfjrWIToFv9WOpLjvKSyraL5Iv8Dk8qEstJYSZWGB+S0P
uY+L0OAgONZV2FOA0VqgujEEleA6sRdmEdmcWE+k+8AF7jhhJIFpkADVMDkQNpvw
lSkDz9t0/8qpbSn6m5UUJvOgR8xlUPyQ6gXqsYigpDA8utRDOc7pOffXH3JBZ/6H
u1/TMMDkLk0c1aontQZqy309ZiMu7REcRu7gev5uKvtnJHlinvAixyVlHb37S6hu
4hprmBOIlRhUZrd5JvbGRv8/o5oHyVx3vjuc9crAttYFTJG+61Q3EFkdeSuAFbq2
BrtSn3oCQCWPbF1z2SoaN8ft+UNPuzCYcPyskWxwOO9byaVDFYmAworpKY326qwB
rLCnIna+ZYLa4A40E+O53W04t2cdA/3hPlWeqcrxGKH9elFsB51xDhokL4G+PwWh
RUtixTgwumVEhxYT8mloQXhsB/XgVIhECiACd/o2zEWfzPb1+BoDa5DudTufZZ1u
iDqjuaNUxXNRaAcisFnidjOOuVKzIjs+kv2nZAaVNpvRjR7jLPT6a6Zubnvnanvz
pAxcZ64ynwowOIP9VQEUFbSg2UdipAsPFgdogloJtPQJbyXeSm7BGw11y4G6zj3H
GNp0RW1UfpPCTJqRcpv9BfQiDDPhBf0WR9xSOLXA3pDfpXnfVwP4CKbf7/+4X5ee
js1tZJh43U8qMHsdFMpbZq5gjFwHOSnllNOEj+HKVGmqJx1PK2jRnuwWqdQCZzfJ
rRi1qCqPJhgFrDGRwrgRwSN3UIW4iETcWE5ArqDQE+c5NCfDtBREnnEJ0OTbyq40
W4t/xNFWmlxB+0RBzf20e3Szf+SbjHOXsj5a4v0YE3YM8gRuCMCzNJdT/dMRQjWN
Ae5lY2MRhP05LFmttOfuXy6rGXxeuxJYXM0tLfl056McucciBpejGIWpRTjsjLzn
BnSihi+3ytaTcJj9ZoSCSQsFSb1jRK/9zcbWCsu+7CvXgcoE9JVneU0CiejHLRiO
SV6NI9wqzI4MEaocFS4G62tui/jeO8d6sxsUb8OpMEfcv5qf8g59GgpAZ8J68J7d
z8vedgyZjRCguy3xeTbvQvx/x/s3XQqgC6d8MFdEkm3XoCZT3DtLyeS6F7HylVYe
bTT1/X8vl0TNQLn7A8Puqg/eWIjcd+cLGUfFOLbA2dUjtDiaFrJeJ+OuyRt9Rao/
0DvZ2Mxk0fA/vKkqzlCyLqsF5e5+emDPtcXQSfwgtx1yo3x05u6yM3nu+SmASooE
gfizlyQ8/CW9jbNK2tluC6piX13Z4GAfIFOqfsc2MANbZ2QngnN7ldLYt/5430r9
20vAnkOf6RlUPEa4TCekThYmxBxCQritCkVcF4Nfn5KZdaFkLc52HVwm29Ls6DSa
iwEH8HoHboKKM2+QS2jB3X7RZQA3oOg7gwxeUSHPmBs7ObUV+FXBzRDbAw0hGL0j
6/bHHcXDCICQKFjW+EYBuTAbkH3GccMGLZpbHrE+28Ltuy5LwyjRqljZwYuA2Jxc
wirj0SA+IoQ7Cy/PHZ9omfaqWeDgV/9Kwdu/A65jAf03t72GRbi9EaQNXPDdDER/
zPq6sCl7x/kjnduVykex6DBTJRiDj1z2F7zETo+/zPRbqV8mCmd13T45PqnX+Sjt
dVylxwqFaBnmP3i/j7JBo/laAxik+vj9RbXVT2NvNxrX1l7/9T2e39SEW0ign9uf
Mk/VN4DepNl3t1wCnNzLHaCOwyIBEGILNmHB8agvsr0bCfVwww6uD8V4MYyW+lie
6dfpNg9m6HUP7XhE0M2vFNgHWxefkq/uGPMWEwuhS/ExkayWHf7Avn/agcAL9xko
8UBcy+VOLp9KIAa++l6v5XQJT2aXYx/M91lu7xWET+0JdxJboE0Wx62L7XScIHFb
DxuhJ7kxfieTn1MKLFo9U+xAOkKG8In3wbRbYBZ1yuE7kfCP4a24qbYXMQdQGzNv
r5+y/+IxignoHbP5gdT0mGVit4jRSMMux4o9+mltmUYcz7q5HypMsd0BzpqIkFD7
lvDxGodxO6STt+2khS61mrzb4IpD1842VoOfkwJtfkXnrs7W5NTU8JFo2/Wr2CJA
bzm7uqtArGWBKZXYYncq24co/vbuX+JzEpXwFi1pEeRxtnThCtraMyGtjiTC/poE
xa+tJaeKyHMNGr9bCFRvgfB/0nZxE2fu8lTHD7sqaXuxX7EOOmoOwYRWbV6LR8ZY
6GrK7ycMNjmx++WXHn4B9d5IHDiKmNfN5ZUK4H7e3mRPhlm53PsU63vWJfRBLQxn
zyhVJX+pdyRrYLqgvUJ+MKBcNYd4xNW+yZ/vRmkZLdVPipz4zMlNrgEjCJbLqA25
nhOkp4TAQeC20ujCsBPQPo3JsDSJQtxU7P0vfxVFSLYSeFt3D2ZTvOQEL8T96p9C
22zPQNUOeqQ7hhxhVRM/qMQ9hixRzcXzJaATIQT5a7TY6IYMH0CaskLUDSkUkeF1
8gp2OyahhgqLWpZaihLJAz4FZr0IqGjFWMHQ5LjTG5hVcq7mRMAEHZFrqmIYKekh
tO3aNsXvVMWK6pptlZSBxv6yH9RAQnkndp+qNtp+AqJui8jS7lAQp9XkdSQB7VnU
dQVmQNcVtrKpX3jEToAX88mQ387sCo0rHqIt6+IzasN424DZVcN1GODRyaurleoH
0ekV5HWcN/wJ3TXOlQnvSCU8qag/L0vjZkY04ZDCIAMO7EZQFbC6ORQmScjazrE9
QulE3nFAwBsJn43hly0AcfDYgJ/ctYZM5Bzavqdw20l6Gv2SOhdFuJZY4sxvI9/i
KwbjBMgQkWTiN8EbzQyxhR+5A+gpYkQn2fSGogCzWYwiBXIV24FeEw/52QvcJXsY
ctpMxfyrifayiJRTKmzGam3426FtfiXtL6DKL557m7f1AzDytD3pU9iW9ZTmff36
7FJmNQIqyPQQpGczS9/2Qj9w7nosiNqqZFsadd8l1mu5fneja9Chgm2f/nWDn6OW
5hxohpv82tJcUgMXkDAEqmIFf7/5TldTJ36LOIjL7vVx7FJgWFqDkHa9na6J6m3d
SxNiJRuAJpYodqgkdY4s/yF0pvP70gHwn3IzoG+G5SOGCkQ2m5FEFcCtSdNjBaf1
p293321vL+94+KiNfZqOYjGVaVLAvsg9ZTItZNrqV4QQTHmV2P9mIkfSOZ61TKfp
WFuqxx/EAKVfrlAck8NbWsz9RZGcndU/UDHBl8bW4NgSnDV1c1gfj1oPDuCgz+N5
NzTMLwmCG3quTsrYnjTkTtJ5i12osMLT1ObnSdedJI17d4W1rZJfJN3NbNV7yIcZ
xGMI3bGolqP2/hhuhF8OAaa4Z7JS4ck1TJcMLwZ1ukSLj0XwxCjNLpOsCS/ohju7
4yUmYCveWAX4tp2PNrYXccfWi/HKDhb1b5jmjR7QK1sFrxuRmKULi73fB+3FwStE
velxElj9UZop9hUr3JP+bevc3uPaqZZ0MXbq8JCTWtZ6i0Vwsp/Y1swlwpDRhSA2
HKaUhzzv3whVjlfmO8arFREaUb5hwuk4i8F1ivULCgzXJSK0UHScdGcoBpE05CQj
Ibal6fQ35XfBvGjPRlFkEZXpBv3UeJlGDoiRQTZhK1a6AcAlK5vyuPB8XynI0m4M
YjAB3kg9ArHveGdsXznd8mKt7kDduyCdzmSn6EazC4PTPSUlRjHh2nEMLMDU6GbJ
OcOftsG/t/S8T2/Pz+9Hp8Zd01SyLQLgIACtprA8Kxu715EK+MPXIZd4963u4iT0
X5qjutwjKnrbGi6y8C1F2VxPmCXmYdpq5aO5WL7RNYYfvdH3J3jrQITPFje5TJQ5
NWYZ0ALW9zAHWCxyvDLkcHIz4X/KKh4gWRV3711Q8uE7OHVe1cZnafdifd1P7ONm
XJRxDFacJoEn6kUGrOtPj2L1Om19rAw55umtHIHTmp1Imi1p8PXHEuRFy1W0y6wS
TQPl8VDVEcwL/OcZnvS0HueogzMPfzwcWVtnto+B9lfxzOUuYPsEeCLF2eLnxOV9
XcNnWlWpf/ImRxwr78MoeqeIQGnaaOeFcsvguIBZsxTA3zWkauuegu35PnNB3mH/
xlNc94EfeZpgzSSN1UnSXdUhXkbMOGMcdMG7yGVLVdd8RgKXV/n6k6WSUrxNXqsp
mP56bq+M6CZ3gCLwE3F1qLM0N0xoLancDEwRL+bfhqVORRcZrD1xYIDhnjs44HBG
56vUm2NXzbzYYKiX8A1S5V+hfLvTWy4rVq/J12390qQ7/q4JAO+cSF/wafmb46I1
oZHdXKPlSetwZq8UjfhBq1QG/VYqC4iYSwv3/vo7YyXMKjugnsT8lZV79yv6H+f7
0EibOAaxGCi7YBQX7Cnuus1jqzJ6ntNjS7jLSPdAdGXda5fDW8mJZczAQ/s7oUnd
75WIpuyrqeNoW0OFEjv+oy34Z258aOC8hHZOjhy8eUspYek4ST39xJzYCKjn8MrH
yxHIeFlK73Ght7Qg8uEKKF2A3VyHi0/eCmAvy8wdq573x9oUD1w1xDo2l7WO44M0
YO9w1gFKgIHaUIBTG72w92YWldbFom9WaVMTQLSE6nwvrz81UmlWduSF6kwpmVnF
eQauxSGsPAZ7AjFuufH2NrSE8Ej518NGOXraOlb8KSy4YU4CuBrib+goFQpgTp5K
yGSFpHBAVLX/DxnDANl72PUeP6q6bBcXdCz2WvhdYe3xrlvkm+7srKVT4XnHnbWU
0MWQFd7IlnKvUlJ/bAmZmNuUfG6SDN752fJGq4+eHQP3I0q7F7Lm8H6OLV8/XDBq
Bc/1Hps72BbMVJF6NI/9Ri3AXY8yA92n+8gQg05wGWR2VHQMyc9Xf1vmC+vC4wTN
D/1C4jBYjYUBMGVuYffadBNqDxOsp0qthyPdYaPUZ3O0rPeeCEkfIm0kDbTPfQ9C
FiWVhIVUpUQeHrJsScQEh8aavs5EBYVc03Cnsi3zCblCitK1Vge2/KHHW2oyYzV3
zyAotNBuGQ0A85sYUzXjRgieHdUpMFAE7cNuVFKorOTDkIwSWVGqTod/xHnLmAi6
vcmT39ERueKBXObhKw8rpbIHZM1+NPYJUcq1TmSfo1mxyj9jqtcvLdeTOuG3eei7
P7V9osjYJl2gytnzakkYDfVaXucyC4ncBCA4roFlMioi0+9Q73ylW0GfK81QOzD2
D4W52F7gZjfJTq5Y3SkpxRL9om199JMnt/ppFZB1GLAlMW8f0G0YGdSp9b5MctEQ
a2IZ65yv1re1qjgnlgDp6V9HR6REtihsKSlzaYeadQNdQbkI0lfWdo4II5k2vU2D
uFQxRKk/CjGY9b66tv314nHBI9fNKCCpprgl5XnsdOUSZ99TuwGIQ2o85CDnF8g1
3CztIBaqUauMrdscuMtd6jJ1PEFxBiRUCy8wUeD1NUIjaXBDtuCoBNA+ytSUO+YZ
mpb2NR6iQ+aocaqz3tdl6whY52gNtnC2XNbTiUerx+XWsIb1GHMw1h4ewIbzNqdM
Ey1y8l/JEFYnJ5TgoldnIX8YPOxCd1fnF8x8Mje346pNZ8Tdl6BVFzZIdTRngMNi
HKlfC5BkTjyRUy1R4DHPk087keovTjeD+GIDeA4yGrGUNOPlNSoNETYv6SZBt1ns
CdWiUqZyMOHDLSpeh/fkTqVPzY/6WZFtpBrvkIkAQbvMl01PIWcUS3jF1fqCQNir
kTd8xOTQi8zY0UGH0hFVG6jejAcSuBLgCC90ONLz2SFmULkssna476CAppbHsqps
OGYrmyg/HDY9KeWGlHzjMylP7Z7uY+rbT4SLWDDN64+0GonHEUITyj1CIMftPy1V
UOJeqrFQ9uS0jF5iAb6HrUn4anKynJH8I9d5SW39OeZ4HXWfPpilq9bt46tU66qX
XaAvOfLzdfMBiNdBD4jEPsmjZcKPcO/ws8Ra4CZegGpYuyLOGdIxNpun8iVfcTxp
7Ca6peN55626EM1E4ll4CP47Pnv6Ux8ggquybjdMUCq8y5qsT9a60ppexaLp6dbl
ZrJxUP8eh4kgWZlyiqNe7ujsoncXDMT58O6njIDBzjDdy9DFoU8fTYcVRcEfRmI/
Jv+hJzIQ7I8rTXQL7Swdmt1a5NOpcSxRR2LYozFhcNMQlzcGYvvahGzJlVtIN2Ff
IfeiR1hUZp3BIQpvpHvqAJ+hZD6eHMhc1zvkPNWp0OCf9GEo4Z6RkdjzLMvZ9bl5
JsKZ/++P/7tIxrPAr2TKQRIhNPIWNiB5k9JP78TzktAKb2UWgUXM+LRus3hDYXFA
PSTSkechk948rusLHPfxosuMc/iDcOCwERmu51fD+ewr1bqd/XcLUjXnXOrdhUMx
aGfgTIYFuT4jwTCzzDkzjaN/Rhs2gQVDgiqUCEQqsnYu/lCW4Po9RnCc8vJMA/7o
xzES81XHmZJGS/sJAggWHIHJNjiuqEWV7yhqSzWdZi8DKGpLjdtg8fZxdl98m9PS
9OhvJr+vqxm7j6pmfGcI/dFmdGohj9sQu0H8ZWPWVB1NnV3zuGn5sQKbpfP6Cs5g
2UtAr/UhaZ/9V3VgW5r3PXqdCnWH5FMNAZ3IGtKwirUKE2BTS635o13BpB670K4Y
HrrDEmyQ//pCRqr3BwZwBfID2IDLZuCznu7PMbg2DQiA0Uio9XGmCEi3KoQU626N
g9UdR1I9Qpm2M54nqvBACVpUvfCCCF/rIRw9A3DDge7325IEcI22wlFifJUURA/4
0kIyeTrrt5tTtBeZp24xDArUd/7N/1wSnC/hB3kcjByPN36dIFh6p2136s5Fidsq
BcSP+JAvNtFSMzWCPnLMoWoxANwUmw9VEEukNrz72gjOoPg1OIN8rRG8BcupTdRn
jCX3bbeqcG8fMkV3mt24MtCoRUqADWl7E8rf4NlqY6cVW3o5gteN5a7A1oIwIAbD
W6T8gwoR9wibPuPWCNuiov9AgyB8KuBwHS8Bb7jdhza5UzmoEbxZL2hrAaP20bty
96wCVYpilT92LH70RROddWEZn6dZb74RDegf2ACQ+2fAG2e/RUGeMAybg8+oNxsG
H/HnGLNMW0+HfgadKYx61E1ghkaJjNPKuT4JSVMn/w/VAaHp0Qc9vmw9eWNpgKCm
6kt/QYm7vJ11BCuAWoQZ+cHFY78Zi7h4svsguRrg4x96latFosMAm8FpmhfvOZBo
QSaN66jSAp8jMaNTy5y1CI/Bpz4FfDOMdEJ2BTgei+9LRNu5VAgLNSu1QhCPIF2F
3yK5rzYA2Pvrd/P/3HwlkCvFH09gpeKsAUv7UsSiL5XUCOgrQuRXb4gNhSrXi7yq
zlynA/jB6IhAZNSoLHY0L0A4SWHOedPW9hc8ub3Dh33foYCzebZeBVSc6tXnLpsh
izv+gUH720uhbDyxqRiFI9aT7xqllUtSRDfaRYxspBL5rlet1om4OmyFHiJFZ5RH
QGgYk7gPsTW+Dy02yQh3d1tnRWrUHNMyaBtIi6DeG0YBOWeA8NiS7DIl4BNbIHrV
//hqzXzZ+UGU42EEh44v4Q0MWPgQ8ZRCDBvnjh95j++VU8qISq+31jq60FsD00ih
KvQagCB4k3L9QW6A7WNQ2u/yR3Pz0h70coCepg8e2r5zicmj3axmvxYC6bIsOW6T
JO6br1Q9C+E+6UP0Pl2BJJLdUfucD3z8MCLQSZb9neRagf3tKSpWAnq4GNNBVcsk
fLUr0o2NcpuQSTt8AOPdWK+rulz1kWiyK7uMqXsvAsKGJ8YI2K9AmbdsNgqPeQ/W
q1a8m3JjujmTGWcu8tr8iDmUJI6ccMxS4CYcNKbIiM+nKyolcSJDgHygMPt088rh
kZ7E7Zq+1kMAVm9IoRfDye5BmiHIwcJuR3qqDOOrhUCbd9XhwU2Z0P9mZCYELmHD
304DJzYjYFyDXzicdWuTEmgwybQY/YihPCbFQizb94YnTO/eO+NCAv1JdPNgK5qV
Xrd6ZIYtC9vhf36cU1/rTPUFLakioikuHwny1uX2JooOYdvsnTJOd9LGdaHanXd6
XYE7uL8i6fLqYQjjql6iD9Rimdpxh4rYogknaCFjDS1UvXsM1BIYrv4TsDSdw7Bl
MOzitw3+LGo8BWnkchhNVQwuQ4GpGMwEHZRe45EwPm9CZabgCa6kk1m1PjRD4+Sv
xosqwHjf4E8slsvASE2XZ7/ZBywkx11E+IHsuOdZUdgCyyGtPN6q/UuBqxUb2CYy
DuBV+PvXauze+Q/2eBLHnUiZYpU204qTm1Q8cWhqv4eQxEVxVQuPtSKRaEh2pMg8
gMqkVLbkStH1rJPxq3Lj3CPpRuds89ZP8q8mopZmObOJ6roi8ivvlNlq3wkXV+OI
rA3BBejORG5+zvB/DX/0GmGMwmG5t4MgawOgU8WThvG0cMxArk/T5UkeR3zD3JT4
ihcmdZDEcNU/1K/CB8jw2KcKrdYPkWYcGVT3evs6Adq0PT6OpmeKmmKvezNVffVF
trzPrfqHAQ0E3AnB5laGyAXtpFZNMNXCJjkr/QC0uw34AhEYhVMSg7OCkxojJBq/
KZgR4ypsvO9oj3syVSwSD2Txgh+3/4dgozESDViJSehpVjnUiemQKsgDY0HWHMkL
8IdcPvR65zXjrRvMpnEazxuouI/5d4TNpjCY9I68fFFegGA+XQKstuFqn+ZXsRCC
vVajtg1Sm2UWH4xD7zTQn9zR7BzrjeUtimPcnUxSz0LPgrciHFj6Z3vGoDLaFkWP
otc+q7mPm/NYVfNg4QhLx+LP1bp3eQVFJKHexJWM3F9YoLqb2TUPUXwT8UqlCVv9
eO4oa2sR+H7bgm0++vDkoe3wyuRBpTg294Esm+NnyZtEisIopSoMjN6M5YDI5axZ
6vEoqpm2mjAej0cxxQiqlnGLa5MfnioSIb0NiLxC7DE5lmUFLFFLlZBZhfIb7eS+
v0It8YjV8PwT97llb1fiW8lVQaYakxMhKNEgPno85P/ZdbizkbZemmCbysQBTusf
pPJv0Ly/ue3RPwwcMEjcfQhjG3FY6CqZHPslgXVqEagZel3qLkAmlq58WyBF2E5p
BhVo50/2BCjuBJNjQbPyOds8TG9IZxI/GPFln0refNHptaNJFafgG27Q/DBIV0B+
gVFYIIGZk6VQFsOE3d1qpe5YrlVA8bJEHO07C7YN9F3d1OKu5yP/JWoqqNUK8c9K
oCO+NTwjv8u2EpM5Zn1kmykGV8lNlGuZXZ8h/5iXpsbWiGjWfB8Hh7osuYjNKHpM
6NE6pX8gJrKfIMntQrX2gODvbRUysNR+3kXxZyS87qfygavtAoEP8QDsDySH1OHa
9B6mawMlJxqB0Z+Id8sUgyxhY8uVLHOooEGdNa3M2wx8D5ofd5zkLC57jAo3ikuw
nq9Urv434SRLCC7QgtOvY0sP/TGW2MGz8NbIxGfWKa+fgLs/InLopVjjmjF0yNLw
YaFISO691eu2NkTzhGuZ0wF0aDfjv/EYb6PoLr+cen03U6hGfJ4UaWRXDWGqSpPi
N8iLdfH1gbkfVPBacmSmeoOP6R7ySkKnjBwrRU2nMhYvvzeGWDXp/y2i4ooaW9L+
fsybmaJvkTWD9P06uOhKflbG3sAaeuC61YcbrvSex5c/I7BqG7iY2tt4C7M8WcQk
1wta+RFMC+XcvRHKAJMTunFYH5dZFRiudNegC6W7qA8nwDPM1DK2pn9KYZOFqXy+
7UF5ch9WZdDSFZVs6wdFrxyqWkmNoO+ol1qTy3AiXN1UKNRpKWIyo0aS1ZLnp6dH
KtuDUMbj7JoGVWDDU0uzJ9JYx847NMmVnOHaMW8jLdnGI1FDxI3oPV2bNEUZ4fpK
CtxwD5yhX3h2ayc3uMj0uFYcW0lfVlYhVenDo6Mp9kgflijaW707GaRm3CDKnotO
SPyNie1R+7rcXGrF3qfdG0XyguGfaTAr7wnyy0B/9w7rBxGbAO8QW8m2iX73qxVc
4rg0Iz/eTop6P3KUCPn8/V6tZDKSRyxpmREBFfMhxLXZbGgBeA7db0navqKELjkv
TAAUYqgNeAnM6u8iCvVAIQUgAb3oD3Z4W0Ij+VuGMJ65xHAryMHN1GZxLXcWtk6Q
rf+TBtTP87O9O0MbWpKad+QJ4TiSTWyO8CAhygucXzfqlRAIZlz2jRdiw/ZMlBo9
Eiu3EMqgy9ChsaOq3lHreDO5sjAcnRNLhCgyjUirWn20OJT9cxIanCl3qA+vbNVm
ukICzNQmZPLXrejjeqOyRiHPJz3++BU5ybzjfuJ0qzM36ZZ4o/uwNKaqoZs96szh
EATsFmSSPIe2IA3s6j5z1dCxw9+98JzV5/V31j0OLFRRHd32Yjt4mKv79hMu6MDi
ApwwgIcK0ZGYwlXokDxLKjWyFd6DpxA/pjQ7bYTHhjEl6/ORxgo/rbyORZ7/nmDv
PXvGf9/Ka75oxw3CWg2K2icQmmEVJ6SDW5qG8sK0aYQquSD2ZefLY7zLo4AphXWS
m9slMYEWTOtmaVyvjozgRdZFrxtUTWwlNWv8BiNpHabMFuE4Jkek6sDoW9BIBM8K
EpOCQz0+wwIUdJHdgkn8hjF7XzLPT09bS75Yl31WsHA5oedMD1GHhaKy0NjdZemU
eN/5sUJb8080eFovkLgnJ5rsxcSKBEn2kaJHsDpPUmUx/+8174whYMJWgV2Nu5Mo
xnGIPo9jSD0X2ZdZa8YjK33zccTg1twt/SWuRqc4TVFPGLsWHxhotEzsVkq2Bgaw
8JXwkePt8qRQ7ZZh1gZsdW0jvRAUNUgw06HobJheSs6Gt24Uo6L4KRkgt8eY+2t0
x3YhdTeU2BgT98Jbn1bZMVTwtKKw4TaskMLC7uvHNLj20HKSbKJaA0tBBRaKjef6
M1PYeOpDjFfk2UQIdMkR4xtLqQrqjW/B878B7KWdUPRYEwSUkE2yxz2XitGMuWMc
tFfmY3vClsBJIahuWEZ5ssBzqI55VlqNm8ipcSXEByuXJwz4BchjvgkNtPrTq8MS
ztJIjd/DVAHLaL8xI5Z1J0KMyfxbV2DySz0IirQqGR9JqJ7vRROZT86k4VVJRnoX
gqrrz5HOt/BcYaZsu/uOvaVkWucq9tDzawuaYIcfE5fmY73Uh2g92+jR9avvO1L9
t33kwdgQYpukIq+33ezDAihSwTfmzvOkH9nEzRD2sTZEi+3a4R/qDtCSgj7KECZC
R/+3moRba3KlyKp+Lj7H4uwhL4oPPzYFPwKfgMk/7uI1Ggi9bsMAotHsRxxuPMZh
KjuPPfNJXe3UexUwfU2BL/za87yWqwyp6wtqiN7kD7/3pooew0q8n1nc7nGzb0pz
6ITOyLL9V/IVPCQwNo8XwLdps3Plw3GFAFT/HtoGWvE1SrWyuuL4P9KKrOIn6fd1
l8EAEGCvEpgXdHFB9oF/uDEfSGpRnkBRsY1U52poLZTnSVENzrsanM4pVx4PXUk1
Pvme2foAJye5y6WSs1ruXFzUgaiWKwxgbqppk7xMikghx0z0XcuNvIULTKtNgqjs
0rwuJUCwikhrfCOAWu/iSp9Y7YpY2Fqt0Gc6p+mPG5I+MAyX8Z1u/3TfHtdPGqrJ
pRJuTnCAbaETPPTSYsB67jE77kTn5T0R+x86elR78t3/BN6NDjtOIgXvE+cjCxbI
qUieUyDqYATVXyvmlGMJgq6MygAaZsP7GC3DKK85zc4FLbsZPK6whVEFU92PG1q5
tMD9p4y8l/OgsZnZQsuVrsf4eYlbxIPcreHZSqQy4wBe6Qso8SfVOJUbg/lhK4AQ
NNEzveg/UpDVfA6IwaBoWR6PFyIjxzVjnn3SROfF/NyGAKn+UpR7xR9ePsxu2vI+
WezfJuhIWWqj1pxmOREUEKlSrDjpA1ggTdhAcNdhJk1GGfr2iOLKyvNvFxCPKTC/
ok5nS05QbD9sIX4j/YF+FrrAZEB47hDRkMU5x2J21F09yYU5LuSIIXJJmnYQAKh6
wow+KIyD0d6AXtKAPjX2U2Wou1TWCVIYvBPEyezqVcU0Mvd50frKmF9QQ5g3pmyj
sSxfKFDeLkyVnRVA93rb+n+qyz0VLlLs931bybcpb60bCa7EwE7TVhA6iOFMZwfy
sYuTbChv6SB81jJDa2LSKfSQStnQ8F/bK2o7Wg5szP20ALpkR5AXKhY5gBd92/ph
XcOsM0SDnYzpllDh/VX/hvBuSeJeXxAIULAQEI6Sojiragq/TFJ829rGujyBzNyq
tjHzPZ0GFcZKbIHplPG53BPMTaPaFVV3qtvy672XYXSCsdWHK14xe41irir5bSP/
3kPIK29S1qClLLT5v+qS4+oKkRJPdqkwttVq7+dqK8atIWxpABT4kHClu3JSslD2
LmuBFkCoUqlLBYPwDTTLBjyreMDPOFUIYuIXP18ZgRC7yNUy3oE+GKFo8fUf5S0r
rMIT7KjHOoDTS3n9eag0NORMKt3ZaTsbCufMrRApNm4HDTyb+npELGIKdCk4hxqN
M/ubtFKE1/5xhnIq1T/qx1jWqR9mN4/pAcZ6apNtTfHj9Ufvh1rNvMnSLz54vjbL
l5nztMVnT/CDudeBDt26ozmC8T7BgL/HQjo4oj82h9cky+iTEbhU1b03KexRmiGY
LI3/eVd/mBV4K2JbkYO4EUqd3AKohI0hYBh1Psm1MkN+u3PBsB8vNdbHxcCfpxkS
W5OXOJvPtb0nsFqe7zEUflByfI/VHlQsWUt45Mu26o56u36vz28KdkoX/+eyM27H
XVek+yQt7lMlr/0UIlXTu9SJe0inv973tF0/VwU65G84uY4wltisG9UVu1RI5OJN
7mk91BHPt9U0jcnU0e2erYM5uaAkRE7m4RrgbplNMOtDbwVfIbhiaZZnKxcW0ZAV
T++FeFCYFo8DTr6Y06R/nKEYYDce8H+5ZzAN0fm3m3x/bX8DM5deeCajw9mGB7ZU
XW+9dq/+a64Qm4BhSTcLBbdQqFZVYGaskJKYOfpLGJuBYfayhRkY+UkBtex4WtKM
Oa3ySjaqUTTIbEDEIUVMfzN9i0KtCJQqeu+t0NJ9qHGur8lt5l1DyCvehOPMVL5c
x8bZ290gP7Tob5FSz+BPdKv4JmAELxh4lLmnULFLzrwRCd1/KY3r3QCbTCJBI+6c
L8hNvSzkYVva9frx5gBkdHyzUGDXfapHVw4SqZQuL3UV58hXnuDwvKj5E2r/lNzB
CsNzAPDS5z5ulEVlQLw5Hud28ny2+knLt0iZ+0hfHHIRy4UWx1JIZhIf2+5RxfqI
73Y0xeUuN62FQPjnMborQlDhl8ARRJRPj6o2B/o5Cq+qUzxMRseos6gZz4UR36W0
yRDleyY5PP3fpzJjjcTU+X8CO2U7rOEA6B8QKyrx+7Vh7HAEXhfRKBRUsc0oKgCh
JtbkZQPdJO+fKLG6Rw0xcn+zyCfiC/EhapGpZwgY4LJxLAu5AldOU2hTg60etjep
SSBcSPlvWe+KvqYKRUYfQMGjmie9X28FwnHV2uXJKxxgfVeoSLn88cszF5PBxIMq
cbPrx12uNX6OhVGQAVRt1bB3rhIA4o34ftcboaL1SxoZ0syRU7SGKYbPZBuDCTEV
ULmKcU3dSCKbLD8W/Ut5NFUr6QhmI1BKHxeihiv56xhTADKHj0jpGor3v4f21EpD
L4IlRdR0ypozU1yFzf9dh1q6+XbsOG1tUHkdJrAY7dRCTqMMp98DklhG9busr/nA
JK6ZVJZ1AggBmHAxMP5Q7iAK5JRTmI4iSZ/2mZICzKadsuWSEcAZTUMnfbrJGoHt
Tr/rVLa+dHDR4P9GaM3JY0X1FCo88vRPJXHvjlZmCbELQB3XJ6oqjezj4cZvYV2p
09XNv5yNWEm2C+OrB4IzaKwov/U8Fi85a2UPdFnRYJyVvxlAch6bJocscx9KpKs7
l1x7XAajhmJPczjQVvc3mpldR8LVMudH/RXNBGBRV0LYoyayzVsBPz+9lrIfJiyh
mNQGCJB5esPkhe75VZqFFxGebbUzOGYAmrTwPaofoRsToLJb9cDPc5J3hU7hCtTh
YjcX27j8G3d9iejUeZ1bWlM/smq7h5is7HwfErrRu5wI3UbaCiPAWjD+n+5iQvpV
e0E6Af+kjVtaz9u6gUyElKs/i4gQfFIPmK31hCLGjzlqteO4/wEazxQggglst3jb
ZaSlKn+zoSnmHUvljFBTb5fIPQNeo8jGCv8TgE13L/AsgQvlSCrHP8f6va7EoB5D
SIzBO34+2ZHHPfYhtbeFS28pkFwi89682/Bk90SP6anRw6v2ZWpaIhoUQWJO65DI
XrlbQiME6hmDWWDbmRjlCH86/i587x0COc17/cHvJXBy2CC1WcwLSIB7MUdb+dGp
YmgEkw9zM/0WJdCYo4fsqF14/XfadTbu3Qt91gkR06T5Z1Fy4uqmK6JVhO9L/Bg9
zN3ZujCxQ9xSQ6rBD9L+fOHycknmFfSh12CMDy7g+vuu5rVpEVTiYdhpBNeIzia1
zUefhcOjSdIdtb4v1FLSxQPd5t4fInm7hZaeLmyrNy/D0viGvDVVI9eyriMb/veb
TTvNHBDYe7TxWd5QLkpuSyBC7nmBPH5dMxxwfY383WanJ0OFprHYvL6K5iGpk6s5
bRJ2Vb3sgKC9QeaXWhKeKesVI4iOJAbV/Uv2ckRBdj2aDK+f16qvYbZENEHiOBzY
6TS59GY7xo7gbkjIwJgJ8R5iup3OHMcwLSMF9k+f4XuGYk7Th9lIhAsiCh9vhsQe
+MCYq9Tm9ncndzQacVPZpwyzFBYiUTxlYTTDVIxF1TXbqE1JJnhVuNyqvzUIIpsb
zUPRpRp+7dXPpdiZllKNO9VHv1Smf7FX+dpxAE6o4uMQsgec3daOHGMYVtgpu7u0
Ggx52Ef5Ja+2kO7ZKXzvJ+fsgxJyNCmRFlk4yCW9EY3VijLdNVBdT1IlMuJcag6l
Nn3zWhNab0aGacUdacUXV+cAEtGhvEvPwpfCuq3UAqW40c+dSl2dmr28R2xbckAE
t8W35COVCTXyn0ogdTmi/gPSwn8xauXd6FwVJgk76PsJ7gePYDKsWBlM6tHc6Grk
A5AWTpHAkvdZtGp2fLfEqLkPgJkSGGVPX0u+ybZpFePNX1gvD/UHPZf3WXnbEPqP
o+nwkP+xYimcrpYuEuGhBIx+LgBDAUGe6WYG+Ro7wUG1/IeIrJgvcDBdCUlZYO1w
m/+CuyMUmapKV65GDWAjCVeHOm51zxN+8N4YsEd9IG6KCc+LMhD7bVsGHfop2OoC
foJcDrRFAbw7UYS+eUkOdEZLFfakS2VAQKf9cOHlK1EztkwLg2oVwcA65I9adqjs
HPUd4uDWgjQAa08SeO1brc/a0h/97sX/bw6nbSnZcdHTo7vMBR5Dn2QO76lidIYE
q8jvAptUCvmsGB1IrI3ZGMwkuVfbZHPxlwIOTldmt7G3bzH/pGXmnDbgSODxOFvX
9GI5XYs5Q+Wx0XkuRGRkpxOs5/z4B9BRGxdMDtwX/G5qiIbym1dImamTV6GFU8A1
IOrnrlH5pYrnZz7mtr21CCHaPZPIRf2/QGeVGOzGGD7WBmvQDwdlsVxj94MxQ7H7
ZIIxeAXbo8IapueOhluwWca+PQ31QQzhD1dmMHL3scReZoctYLbrqu/7wCIW3A9U
UFgdXES0oVOwLDKnqWXhK9QYagVGbbclTg1dXcxHZyX+U7qyiyWtY+2wfgrfKogP
CXKFZqkQ2XwW0E8ygA/a/dhDCtMJXs04s9VuIyjSwxZC7ZYWRpYlt19dUZMlNbbe
YylQQ+eGz5+B6RCOqXqCj7pJzyEzg9mjB8VvuTsumbtlx2UN6g9lSy5Aiyi2sHVU
G7Dxs6AY5GQ8bQQDvRJGQfvPqvi7ibPWT+IJD9R8GUk6JWWKYYdHrCKSozaQsflx
slAKiotewV9JteMj5fi0T0KG6bMeRDpcWyDr9mxyykC9WD+QmRHMMkLA9BXE8gH5
trlT0hNy0TudZOMmzsAJdYz6fYjiVgLpAvc+p7mZ3EBQZk7s3YeNw8PPoxrCxvT9
R+5BRxrf2BWZ+ne7xlQBx3TlBTfPcvo74lsfp1n2numkMO9dWMtfVzIBng4S4kZd
wDWjNZyBHHLnYRIDw0Igs5Iq+MzJbrYMTmuHv6/qS2uKVZ9Dsl7Xq5SIm/83D2jg
WlJCIhMRkm2cDtB4T/lRVCqhn8JgNNYH3dk4H+wnFN1bH8JfblQ8EqWGp4jFVX5s
/6EMFN1uNpXrZVW/Jq8m+COvTe0phXkdrXeXSR8h3H7G8dBd7PIKmi68IBVuqhkU
1pGFUuV2x4h3BIFUDV1ghiw7KPGLLUbBi2SzRZliFhYcPA2zX0bwHIbeMw6i+VXd
ai3j4/et9f4OWpV7OvPceCVswhzPs8tEo3GWGu6M/WeeejJxHreBPgJKqgOB/BnH
2Ng7vb/TAHGTBQaicXOnhQHhMEimbxga1Y9uFduS8KJXy7Mcgd8CmxcBKsqmetPq
YYoyEmWKyr36An9wnltuWqAlWfbl2y6pkkZe3VUjMr4CmvXfy+EOWK0Ip/12nRE1
OkuwauMC88Ssh2h/vlLrgQGBPZrEjgTJxDhc8DRUSYL7VgTn3wrLNWG7JowdHCcU
jYq78ABMcfXIfX3DCZ0wjH78mX633mO58YcYHhYIn47Wm3Kj3BvCZ0emtJvGd+UV
do7M6XZS0d8I0GfgZJ0VIQP8Q/t+9L8KLJ/LaZT9WSdAEXS7HsscsIyt6EY7SKMU
2dfq5NMSW7VfqkfwEy6MKt0HHNuQRtE6ahXu/8UmZEbdmQKtbfbfgBk4ClM4EyMY
/Te4SjorPS73QGLY/SPHNzpOEZmtacWT1WdMnqHbXMOdBja6M2Xb5/UoczAzFkLq
f9WP03/Ra7ZaLNZ4rRMiqPhdjwv5xP68tlZ54+EYFmfislKsnZD5wSfogkULdw5n
Pzhw6UaeZfyHVJhGRXAuUqERR7mOwxljRmytbjjn0OGqv6GLyEuL998YoCbye0+p
wWJZTqAlZDRott65ut0iJkD/kDjSk6pMdwRyCyoXkRZBmmSv6JldK2SOVtfGVo3c
SoGRmUUmYgSjvjExSNlS48K7dJRyaBnFhF6X94YF9P13aC5NXXwFH4hfPYyRDd7j
mtrhWOE9QH1HlS7zmZRv7K8zOCvApSAL0TJJb9fO6V5mGyGHfinRw6RslZq/JlbA
IggDX67EKQ9CT3m1XyaK2hS3ETG9B74NxpcsFzEuv/WYcKdYRVgeO+EGsewrlF9o
+FZbTPMCRrP3dOk5K9KVRqdVkqkS3iH2+xbXmrYk5SISYS5S+yCD6kpaltMeQply
zMKeZ9S8JcJXWuI7Ev6mDeICvpvm8vwjaGbnZPPFBrod5rrOXgO+aFbvVJMLxNfA
pr0evqkwSfnpMnNB9l5TB3R1/Rx0PmVl/c9O6I5ZQDXrIhQt3lB+IpT+CvaePE3z
g90UM9Gxd+5R/waatBU7SpjOhW5Iq+BGnZmXGBJIha+BnSWy2Tp5DusU/dX8qbp6
sdHY8ZAEPwTlcFHnlvzqJ4pS5UzaL3BNtaVvG6XHqAjwf67u7BgXH5fX/R/KlsNz
F/YNyIePLRyT2mVUxzvwXuZnRulc6z1kM8yKeheewmg7s1ZszbDM7pUQ9ddA/BLV
EnvBqQspxOi22Y+r1KGSuqcKf38WSf0d0myY5cN7zfGg93wSsu5UWwZpLNJT8Tzk
/ZV7h6/N4NUNCHSVeLC79nbHbZnrwnyUXAzZFG7FvWTq4+SKfAXnIAwqCvmWMfpc
mb9q3xFXOBJFj+IumdUDRr9hCHKL/EIxYmaAC+GsSh8kzUqT+dbyJrdi/bDjU7Qn
BjvCV6CvqcSsEo8AvW68l6UrQLCiMiVu1lPnwfsX25wGuvP8dnhODYXp3b2OY9Gp
BHH1SqlROF2XrCkTvhATrdufJCyVFPX0vUYqsJxMb6e5ntSY370pG2Z6cOj1eydO
5wZEsGDUHaMzYUHpQz5xBusp1H5SjQ9xCIwNI5XfHeDE7qtaiDJt8Hbe6z00Bcp/
DyaSfEmCrQjhoBoTSQXKugLiBx1utOEh3bhRYH9R4CB8Us2r//x23LmKffPe+/A1
GjamIe1L37sINZOstSTnZlR2xAmxrKGyv5CZM5oKKCx1WagrzCLwLrbPBcE/IDFN
9GkaNB4ksrSEruUZzQbbihiPgkuY2m3Kkh5afbGKqt6rMV0+fBHoWJUDj4wX2hi3
EX55+L1IfqkxVYD141e3NF1Zmexu5oBoR8H3ZwrlVyItow7Blhr944zLc/XEfBub
jip9Qwi/arfSeiuDmm2OvLMwLTNAgqAEDfQahJybM3n94+u3IaOJPQgS5EuD575+
LdZ3Wx4e9Bta1fZCaFz6fHElvpbMd7eyEYprIA0qWIhEI1xYtM4GPq0etWOF3BES
TkmtZDgUdSRKIwKLsHeGtD8w0OlBOcQ6/RCvI8Sl6JMWqllmpuH89Tq7BU+n8clB
9iCuJezo0SDb67IBs3bD3z9xLmf8sXYRs54a68WbIbXow+fRcEp/FQysW8MDvM2S
OHRGS00lvkUCEsrirZe39KrCw5WeLn6/c99dMc1HhAFmHqAZWE9fDHSFIrYp5kmS
Az961/8TkRjlQjDjwIq13difQvBwM+0Zl/DeGae+EVMo2F2XABXahkNDsfsJ2VvN
1JZ1H7UhXZdYr/W4cQJyiLR/wutCr4CexdgCtBkSLOjGuP4ntQjR5db7pxO7qTkw
HUeKxeNy5f80lbtYkQCj6hAo8/fRasK1N7wWtu5yMS8qZmTswxAk82LvTdih5cZ7
KxL0w9ygOymKhNveVQmLcsXngvqqlq3AtAJoyVfuKp3A3NrNmAn1CgkWiOtlVip9
KIRKnKxsy0RdkUdegQo0UfDUL6jPFEz+88MdjUjc3VW04DKB6YU29F/6uSboDMa4
uSgQRojI6oYiQ3SeklfbFzbIIYF3HK090WNN/Z7ZBRDrTeLscrFGcxvF1z2RYwT7
V75DP3htFu8IRrVka+Gze7JJZWcQwC146GY6OcJRPtjbQTmtM+ElWsfyYAEsxMtu
LhdgoXHSiFA6M2U+Q0W9xjhpRjOFcpkCxijnOmbfHk4SY5es6RZwmAChZcInovJy
3sTPlUFkfT/fZVYJsJkT2k4MFEq0POGnnpy0k7/LkV33JZqezEj+Hzf6JuRoQ0N+
ivW4m56/kIjFHalF2PPX67omcAmy7YJNfWztpDIT7TpPij9j5t69uOcRPhztgOcT
LOKy0yhIL1hPAfDHG4fAFeMZN2sp2qNjAva6BA4CKWwOk2neJJbt+mMg2Qsczotx
dbs5Vd2ePO9StO2PsyT5ixuehNSW+2FG0B6aDTFdzt06wAA63Or56kzNuM+c5yMy
BtbqrzBNmMBqe7KjgKNnBDOj+1+pdA2OKxCt6KUepEnAhc7rkJz1reqZjI4C8BsY
vmVpWjTYqpr1a9snsqAeZA1yL1NW5wAbmITRAKF4D6x7BSPUyr6t6aCix+CIZMH0
lPvuuiziCtnsSZlP+EAx/DS0f7I65Pl0PvEilhOkNZhbP9Ft36mTjt68nm5rVT+v
4nGMjwdLvBJ9eYRTjaaIzYHh2FI2B/yoqA1X2/UGGc4o0+A08SLyIHdjk6m3frzP
+/XEftj+aXnRrHF5KQctconnM0rje/xyNDJ7w9Gw2ghGvLGIqFK3QwL6Gv+rEBhT
OGBvLx3WXbP8qzkXbfoDVKzLosKbVYUTS/LF/TNUDDgoLHWEtidWksvyv/UKigaT
0kawttXziTVZSxZFYRTx4dqV0AqnpIs0lkK56OnDhrKi62akPHBwNH7Xg6BGUqY9
wvptF6fWa36Pv3jZpQAYn4BqxoURXdazKgmRkM4G8w15PzKxt59S10Xfjm8U/4NL
UPQcZ6C01fZaarSvf+VO3TThoolCz1IggEz/vx5r7yig64K8BeUifrQYf+RxphFJ
u0gtze8DCZFCX8sbMFLd0zHZpp3pJnnfXTnIjulUgCnpQgHqzHbOODygi9MWSpaJ
84xJYXPeYlw+jczKn4Qgv7LyYQYLTBmxJeGix/4w7tdm3CI4lx6aqDcGL0jfrzB9
ZJSGKJdWgB/onILij2QyIpBVAE3jPVs5jZgcFtAKyFO7DTEV3JQo4xqA1R0MBFil
TeuUuZ/90xZKHrkUrJKbRfNh4fiqD/5zHPyTJSTPXrn1MtgvAGFQwSXUKmq7wIDp
1QU4V6Op/mqauvowJHhOuzW6mE2UZpp2ztAzXJ2rV/WDQW9z1Urd9aAoJlU2599q
i5Kzsw72jSWyDdF1uKZVjjc7MUFbQJzKq6hsMeuVcq8jeTJ3JdzCgU1lCq1Paen5
lfs28R3z2LUfT5q5XnLac4p86JnpurUeOMP809gFQ38f1Y4dLUIByO00lK9IwklP
3enDmEJF1yWr9SysEFGrU86BuR217gbWN7DxX82HBXx/ep6y05st4GR6q7J/yx7j
QJWJXaog9mSUQntfYT9m3TtIxSSgH5OG5zUtCEKCE3Pgaz6gCT5T8MdXHBu17zYc
GSr93w89OwSvDUjH6F4EB4cNbCJH2VaKjeZBpxZWl32SnUtd5C7UEgBd0lkdvYMy
+QgqeWxgPbqmwooIGFKO3FGy6v/mLN2f3rTEuvhZbarzlqe2zkIGbl0m2YTL92jJ
D36h9EM8B3f4gwz0N7SEidhZtrjIVjmxkz5jVN7dlftacfEdksyT3awJAV+0l/L/
sKUZiPjLjJyLu2ncLtc+1s+D9Clj95kbUZbBMwaN8L/PyHFxayGtaCuarw6yiR2Y
VxPbd9gKhdTwLXOpJPdhfPM2KbMoB0UAKsK18znXpA0ppH+TT9VcW31HHeI/He1G
xVCMz4KeICeEbq5rIuE4auCQzjdi2ptiiNQi9eBHwhlSeujLjUQaAUnEsUtyYGbF
SoeYMkvQNWk3LNpGFZbU/DWdhXx3JraE3yQh1TvHafb8htF8sh5nvpN6oRJY8r+/
YvKOGZnVt1w73OSvhwaVcMZb21k/RDXJ6j1dw9ttugQu2zEyZXejQ5SLvpMPQlBf
5RSNnTiXwvBh0pJuomK8gOCms8yYHr01zv8SPA+y2q1IXQq5ynDo0pwMGAM1+x78
icOBqpfnEilII0qZtp4yxbz1AlP4mAHPQlmXRzL/RI42wOMf+LymmmHGlF//ZlO/
2Z4Ld4YQsO9GWI+qArDnz+4IuNNkm+2SoN4UQOHlYgI3lh7W2kaAJijBCZcs7Vvp
JKl42Ms8tQBIGVqES149N9XZpWN+qSka0JBTkGFbXY2D+gbIcmpIjPmN1CVQGhAf
jMkTfb+7VeRpVcik9nKjJZFNB1+YTT6SiUwH7aEYzHMrJ5ByU7oLSa6oOGSuBxyE
BLHHjlu8/a5U9slse2uc3OFJal8Bm6oPu30oERRt5Q8qxvYMKBPJ5MEiIwxg+9Yh
tQoTpk7lsMtVcWAwND250UVZis3lAAq2ukX9sjjhbnZogWALPf6vJR43tW24Rj7E
8U47GbG4vodmnz5FC7xVsCECTlOMjuTYcPwHbRExHxmH3XjZWTsoY7ef1Jo9O4uk
XN84ma0g+0cdPm/8o+ELTu9el7qtH6/S9tIz4KXmsJCa4Ovoo1l7s+1McNiQ9Ojl
QnVIQLPwK3TsVGU96ORQsA==
//pragma protect end_data_block
//pragma protect digest_block
0EDRWncZMdAj502BDnQW5mm9MYw=
//pragma protect end_digest_block
//pragma protect end_protected
