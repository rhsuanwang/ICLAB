//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
IBTozFAnVKFooqZ2+EBysy91k1ICrJCeXSVPhKsl4gIHWsjAZfzfv/vFnF4GkjJ7
YMECHxUX3QtD0YG9RRDyt1/UbaCvnWsLEKtavjFP1+gClDQJVHfyXdfFSb5uwBIJ
drA1u52pbXLCIUobZYeU1dVE26o/OMiu/WlnO7IPT5UaNdLE/PVKHA==
//pragma protect end_key_block
//pragma protect digest_block
XmWBiOZ8FswnvF9EMCzod0iFtek=
//pragma protect end_digest_block
//pragma protect data_block
idkC39usqhF8MoUUMfmM1+vY4WUvuHPTgNlEhr6eUCTcozDhRDPfdeOIiwSSPELM
3AhZssi3kb5JvgKBB0IxHX6DviW0GZuZe3PAYxQcWvgaELXjLntGiwnBpqEpfVzw
PCNExQMBhLtmtV63t5Y0h71Ll/brvSc25mzF3rUsQaFnWxSaPu6oQe2Qwo99Och9
w5MqeJ6GMbXQ5j1leH8YOtpNcHEL0jIRArvM5T7eWGgJhKGQNyVLi1phKZk1+4hw
qCqOW1O/JndV4AOSx7RPIxPpY/WSsCzLhJiohEio14TPDSQPi49MN+IXQ5geRvU8
j8eT4T//JJMVtcC3yjj0KQ==
//pragma protect end_data_block
//pragma protect digest_block
atTYjHQbhrRrPyb9iWzpIyuoy3A=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3Rwb6r6gcS9PyvMipRPMDXaMGI0ebUdWt/GPMYAwIU2kZy/6IhzNTfYWAxd9mwd4
JC+hvtFQZNtxetITDxQU9FqRol8d+vaUUOYdIM/PYCoanGjzbGr1CqOnr1GrM41e
b1ePFZMVHQ4VHb1VzclG6ZBYF9Vc+IzjWECFXJiyJUnzDUPaCCH1AA==
//pragma protect end_key_block
//pragma protect digest_block
helaAI3lmkPiYiBmJewZCTCD6XU=
//pragma protect end_digest_block
//pragma protect data_block
UfK1ZUp9YoJGL1SvtPEcWkiP5mcTrhorUv9ZYtTaemjP25cBCgqiHKP9T6bA1KPd
0QQHkWXumwwj6HQ/Uqwq0zySUzNR6uOErLfXWa298VjZMLFtnpj9RSIcCXsrRfcG
FCTiRdAFECtPfHXKC/ZJy0O6pGQExoeJw1POWjLTeQM+IQmcI0p3koa1Z2r8b9Nv
w3BZQKZvMntqbbYWUaRR+cLLsDW7A1LeWL7q5ZMCVL232moB2I1EHlrkaMTTOPU2
CmO7Q6WRFVVop2D9wSIt0v/uXBtPo6okzL2IO2fNJdD60UkqiyM0nwG0Hz6sJLYG
HSCeFRkUOCnILnfSaMjjww==
//pragma protect end_data_block
//pragma protect digest_block
pfLziUw9PBeugJogCZ1MoYHleg4=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GB5LgIV1u8GN20wTMc88VIQjyHbkSkvNpnmsd+RMdgOuiBRMA4knh+P4Pa3nN1Yp
h+TOk5/ys3H+HpZPfkB0C43OsSpAyHhNuWJ3NhwWVyt45K5hvDZCPPgvVm6SDSeV
2213J8Ote1qcWbxt4f+NYfBpbi+ElVSRLQstjRJ80WeOOYi31q7xgg==
//pragma protect end_key_block
//pragma protect digest_block
+ICUCwZWy4u+wVhmEgegQ+YRFoo=
//pragma protect end_digest_block
//pragma protect data_block
apKtcohk651+o6aTLaVLY/ZMji2TmHGQzyKzgOa9ey7iuJz5T4gPIxY21aLhRl7w
IhHhXjkxRU9PiQH/tEH9Kgsdg+jqqbHLgGyEo7vd3pDNez5GtF8mI54XJoPdHMYk
rmOR5RTaUrHq0GY9yRpMPHq8a28HQCvIlx9R45N2024mcDfEto2u1EsSH+a4mWyR
r6unuhDYiuW/A/cyjeT3MXiOv4mX99bRbSaXTNMQhRT7BZxjVbeyUbkuq5auQ1dQ
QxvNlyIY+TvLILEPcxXOFpfRonNvO8P+sAyv2O2voEC+AVksGzBaRGlTjuM2x9kZ
O2tbQ1mDLHpEZ1G0NBwPxQymlcQAnsQyw+Ijelab5OuApUtqNaqDg1oBIFXrKUqS
60nmIFqxab80H3YRzg7sLcikriVrDS6SoH7ifL3zesOwfpgrpw9wLgLnpgvl7XBb
X86ifGygTg1V1EVUA0yjzlTpLKOUx6BMPDLMVm6ag0Fppkp26aSUXDIb2HAF7Qlf
CFd1PJ0AR/Oy5aBETyivr++b2f4tAFcaGMoFodKzV5Qce1AMfrpUKozw68c6Z2/i
1zoBFswOiJY48mF0n3IS2pRPYKl4QNfi43m64uIvj4f6KRKJ/kdZqnIHYKpDA65l
TVgAS9t0w3V68CdQuFSOLE0KibEtBClfMJzrlIkBgQXKNi2Pbe8MusQlEc5RmhNS
T0OByV2XnQbzi3Nj5sFeSGEBgqxqyTQS1hztODb5x+BwGmIbNzsSxM0YKk1QNmVs
fIhrATjPODKZAQVRHjISI2vPDS7n/pXoXYMn7jOPCR4I01IBayuhyuRFr9Fx1Iu1
ZkOj7RZEsZ5kLDm6ZwRnKyqChhS7KuR4D6LO/+9fahSGS6V4ixOcbUe4un8D+x9E
ymAjr2Y+l4Xn1J/S0s59GoWlqcqlByMo3MDdcdbgfwTavQ2KvGvaRdTEF/YQsIHU
Q/cFQ+ig8mbr7mXrvzPWQM6jtftDglTznzccezJb4EniuJyW6Pu5tL8w0yCD/60e
NldAlozNOj3dH2fImdKuLi43uiTDWgh8cmLpoq/y7i1VNyKT3JRYV5b40xkhDlWp
lwoixaFHU8bavFNJ4kQ15wN3hxt7p9Z2fAB8/QJrsTebNoOYhc087XqWi2gcWChu
bFNd/75X6ZwgTGcfmLfkdlcQ09k6fixmOIwKIabTXrMjzw4osiktoTqMUn+goYcB
U2Ikewl/rqoEnxabLluyGzG9uVcaAQWOSmgx3+Ac+XS85uwEM+J3SCCkHOMflDlF
RBLs7ZYHyaCepEUAHAKNBfcHyVbQf6EJer7M5sco1NiChlolbbwjRUJa+1A8Lzcj
7IBihUl9Cs0MJnUMC+uBRaLn+r1/HqsJmajZgw4puIAGJaXVeNUVJtEPEDDikJCh
aXMSaTHWmPsyR4SoFTNfv76+o3wZanpV755St2nQwQO5FC4V9NRRAL4l/ZfSdfN3
a8NvbgaL8uQoHNCrAuc4EexqaDoNxx7w+4lKPpgZMigihn9FicC9L1zUpW5td9Gc
OU8TBX3khxUgajOBXJ8Z/leAlkEkhzViYGWURx0iufWk29HGUX5wxSQrekiFTOIj
Rd9oFJ0XfqMKlPCmoV0wScRyJngofpNfqBw1cALyEW3DSWyMQY06mbr3DPe8WzIb
BF5lkhnKZEzy6WHWOkbyBLbSJd/rPhbDgtFkt//ZGtcXMGNj9+8ENWDTk7fLsm50
7b9Pk/wgj28R/QRHuPLV6aKGog4zpCV2K17P9ZaNdWnZrNQHZT3067sdysl83ja6
R2izEE9xpWFnoFjxVhpJvepQMbPd2GZEI8KclTTAxsJQe358iGcX6Q96xvZl4UiL
PNTHuNFNLKyjHVlHKX/AHqeOffKUxIvzAk6hpTKuofGcSrPkxqsVN1GrX7XiQkyY
urH/BC1zYefQw5GOzE8NFdXzjt9nJn43pJMADWdcWbiXwzY8RzlWm3VvUxFzTzOF
1W+y4yahRNeFRSIRVE+LZ6QPzW0NbhiU24KnoT5vaiT1pR+m4rC9D9h2+sA1HOHN
Q2P651k1LrXWgvNJMs4miX8wzaIhT6IrfGLMLJtTSBrm4m3Vz0tUyNArK/fK1o5s
iCduDZXk5JprH9Q73xpqcVdowtr5sLRuOIL1WNPPal6wgq0VplhYbtOPI7NrvCyB
lnA5eKu4dDRDFMqdjU8cnAaQyyGjsJaNDXS+3vhPOYRi3Az7q/2MB0qlq9MyIE97
LlRKcEO+ts9sHyXGCVaxTq+TDa4RUkFYSjA3RCaaV2fbaEtUF4DfCg0vOPwdN7eS
RkhYBTo0sgpvUMuxPtO+roWCpmgp1YVNFStkmTBwL4Ma8WxLjZrTaYuSmQYb/P81
CaPunQCk5Asqc0hTzi9m/K2dUM06ZzgmWcUSAd3S+SR6k995Dmmm1iYfPZg7GPf1
kfF2Msl+FH+w5qDlZ12A/+P0UHKp6rlBmCTgvdYdKX7C2ZxkHSjQC9qTc3NPpmMG
nZP44MRJU1/p+0FBxwH8L5y/Ebq2p5YuUNBLOFDf66tRIWwxiMbrDKIJLamEAu2p
Y8tYPT1MMsbPJacOHVOr4GYJ0BLD1N7FJ5MGcsnLy+v9y+u5aNjYXiQJ5q1WPfr0
x4lR0J2Bg6MnWxMADgdvJ70I92oaB2lvXvIkndUXZdZq9qVoIyvzPsb+t0rxA2LP
bnBBF+hXXXk2OTi+jFCs5vshahW3XLA0Lov900qS5yVyvwQyvyd1pydake8aaZUm
Pn6UHM1nrlsf3diSWTZhWAb99w1Pomx94xiEpyf5Mn1/A4ghEG7GkV6SDF2RsiFl
Q5imGPDZr9XqKbzu9hVWm2Jwc2EPhHEcqA9cYel8ednlho07I3y4cQiZBvXBAuEc
LPztRT+87cV7aCL6DAHOhpyU7UBaI6GwnfP7R4VgrwJwtx49BNsQf8RMyFrkQp3z
QrwFR4pOHqi9GeJV9y6cq4tIhvjHGhaUg8HIflKuEceajhXavOS1Q014BYmnyciG
k8opZuonDdlnmstPDjDWPBohnzvHZhF5WmqONQDJ/fOYU8RiXMFk1CQ9G+gt8bAC
/EElFpSzPUutaPkbdHCn+7OWAVX0oui8tBsnJwik8BVDNVGw4E9xeKhOJLx+p+0y
dEoDEFPxd+NON57VtoMURmtJH6lHkwdosAPMfnfET4xvBZbljgiPuNZuYxF/IPN7
ROZOJf4z40103Kv/tu2qyxQUOHQ0rs2xlVOfjsr0tiaJGv/ue8a5yCbfRElBFA2C
vGyaMAYFqUEtKyHwRU2dv7e7za4cojY+3xf2lwpFZFHjtGAUHSeKQwH8E+gigLTw
8BJadqwzSo/h5hN8FDjgOAJvTbe89leoibBKDtvYMkOHWQpVtm1SqMcvxtSxnsca
i+4V3thm73G2KTP2L0n2Nf/T1I+L5uo2+yMc6YtUpW5TaZqjXvEmNiiA+g0/25Ve
+3iYgVkaj8f/f7R2JyfnlmV+vdWQq5raBRf7KEdJzOoMsghnCL7tJlc4BFpDf3qz
1qRViBEmxIvS2EFb1dKtdMh+LPTc4iOV6mz7uoF3dTTIENG5/aZaNsMdDwPHwJ/d
Y46E2uQ1PGJD7Tq03PG2qPae3B4Vi87WdcCfdQ62CZBVXrkA+fMIPuLKktap1lLc
+fL+P8F3nnuwwjIdAZQ0WAWWiS/41KpgoThwVQORgALJOgiatdoXcynTZJSE2a4R
ERXDm9MZ/lkgMIMM2bVQFfKkctEolQ+B/hijy9oVxN0uoDw+UQeBFNW0GTeOh7xN
AKy1CSKC6C/wraHaOj2wH5KlRGNV+scdn5DjGsWBbNxfotT/l0R6KWqVx4o3ndmC
BcOC9JOAjLffpdFoJsMQSE1YoazKfOUpT2qnBCE5PvRzbCF+cTtbtDoNYL+j/5wj
PwVAuXCTlfoz7uHKQkhuYty9nyOpoTeLgxTvbhp9AdgdTRw/viMTTKCu0+q7y2AG
iMnjgJTIvNTeIBC5Axjja4TzPlNbgMbIu9JT85Pn7QvHZK2egIa0Yr6+Z1L11WRc
RpukiPMmCvN2TAMev9prbSKBrqn30+cua8xsNtZH5Cg83S9b5A36xc5suRK38ZJS
hRzpvRMcfkP1A0wqxYBrUL5jvduLzB5DDPC6+HvFLwTdHCn4DxevhigXA8KaMA2n
Yyu8jjMlqX8hvBisU7RT3UzAAeE8pXlRei4rQjIuABGB5bwuyY9m5Xg2ix717ztH
EciEcWbVrByGGZzRqmKis1SF/YIRmXGn/RQbgiaAwFq3R/EgwNvA0KjDR8/gEIRk
6F8Rl+J5SgDy+AVtYlSMT3x3FILiceCoK2VzQXoG2mr3Un2UNERhymgxfQcJIJvE
/Nr7bQP/Tn3sJHwjjFSU1Ji4mkRZlvo03N1LluA9jMtc22ptPnQwCAtNrR/HIkaq
ycO7GxtsuueBIend/kDG3lbX97B6Kpb1Navbg2SrfvVd+12XWDXie/7+v4kuD34q
Hu49oLPkgX+vuUablrG4ZBe1PP2kTaF9mijw9g8QeCuKQO0fUQmWn1gO5o8P+zM6
yWcxCLiipIcRIBjgo6uM10a+V8OaVlvaukL56FQoCLRdls+SQw0oNSFjDiPqnQzi
1kvenqadNKuekTMVIdb5H4mo8dMBpRPD0qYzD6MxlWsYedce98T6OoG68M2Cucsf
eD2BkvBqiUcEV5V3Z1sv/sReBS0FtF6+plRyVsUpCjhmEvzPJnhiFacBzUBtFLSI
bfEzI9zYnVoCz48idyau21Y2HhfIQdIiUftPM0qBMev3C8CcfYc3dL4dDcoTboCt
Al92gNAgtxKNyMox/3cRxhcGYa42mLSvJTrwEqQkKxpH1EyNOxq53/LyG5hmH+2g
XKsgmOHdEWafBPVBkmndt+KSpZGhXr0UgsxGBjjXImVyRDbZ+4Zm2BNMLal/IYM3
BooY+ehJEobHuu7X3/x2g0u555GztOsD6+14m+GJu+nczwDV9uiF1B9JEhi7+n/F
Nb9vRgEUBn4U6QcZq9k5ZuW+i6d8Iah1obLH34yppud32TaaLpXGO9jSZDWijvYr
jfdTTezeE9kx3pQLu73agrlF4hFOUciM3FSk4zqa1cdWhDeu8gwi+Nw8u0Sw4FUR
jQv3iBqoAw8P+7EwEK1UCYpWKKIGsuQf3JLEOBL2C+0p4hA/qhd4/aj+/WOWTZQZ
9KqltRpeHMmT/jTpOMQm03c3R2tIyc2p9AvIiGH2ucYzExRg4lRRCiL4Uxs4L1Oz
694302oVW3p2zSrbj+mF5E2rlS3LBuaDkW4tPOOyuV0F6JpdMNmSZAJW9X3JsB2l
7oO687UV4F8kAOvzkC2E4L4J70X7mGYXIMOxmdjKbeS7nv7pp67Oo2VXm0rpp5IC
wMBtOq0b/09cmKX9jqosHc8pFTFNcMJ5pJOSLoS7hChfXwDomCX8WQ6jbDo1IA0n
7B/eMS2pBwE78ZzInP3Tut0WO8BLsnN2uHngwqErrVVaq1Cudo2AdeoRmoWHesid
sRVPyCT6FmxgNJnJfh+0uMapISWOurRjIGABqw0yp1UHZsGFK/n3bdokasS9rOud
S3+o09QDX/j42/SduiBlQHswdyDlQpSUUSun43OHjOYzfs5LBJGiSBR84YZkLPTG
5JmO3FaGaZ8F2cJF8ENZNaNh5fSAQFeLEd2UAj+FwU19RWiLD7iis9n4PwdG91tO
WmKSGqPZP4EgdS2MGuWfEpqPcB29MxRawSiwafpyGFhsSVMdCDLvH5htsW/dn2dH
gU0yJh0wqodGBFbz0dbXpnuzKX0EhwypfPS0b8Wyb+NrnAnfvk6LMgPSbkJZS2bw
4cdDn2ssgnTWnrHUS0Q1OAa5pYBA/HUl6FsjoNE1T2rp/ydyrGLV5Gla2vijLQr1
Uzo88qpaxEj1RzAy2JAcONr619J8UiQcwjFUWVYAF2rvcQbKRH+0TOHMMLu8J1s9
fhdN5K3eQdLygYFN6JrpjnvfLYnQAswzxfYuc+OIyHHdI+umL6rVFqIwciBA8ROl
zuMTY6I+yq216mvkrJ3vjaxs25iIWglpTAz9ayuXmNKGpk/I4KwG0+iihwgLFecG
xcwYpvzRwC1TXqi2ZR5DZPH/riES61COJh2Y3/3N7yGdtXItLJSgXe3q5u1+beYn
XWadXOwidrmfvLbTN3DnwCii4CUbWNk9zKy98TLib9cT5EQPDOa+Kfnfi1Ps8T7o
ltQhEmeue5G2yMfx36833L6GvGxzL0GtU9F5i4gdhQQf6UUfvaiSjcyqJYCRBpaN
AIh0Xb7v+2bcwUkOLOzAfVMdCcvQEYQnUTbt5iYx1hB/NGAbFJysmI64gANSRtO/
sATCk3sEILkfOMgjgOzAWawIUlkcrXwm8HR+3AsS6+FNc3VI7oCkfZmOFQJyrR6x
6bbhqtSJSOPMVPP9Sj4LK5DKEqXS7o5eS1BhlJdAEXkZD43Znqu7fKBOR7HFfRqJ
0xLP89cu3aYEB683QsiYkJ0L0zfkJO47aqzehTlqjUbcs+YUUng4Kgv3Uzx3w+4b
nhb4FjwpZ9eoMNuBVMxIyyY4GVlJstEjSymkx45n/sFhD+YXggIdxryeYH2uGVZh
ZxWaIJ8omLzoOwvjbWEW0cAx8y5UUAD/ni5Ok4gOWm2fP7PDyMeig3X22PlUJw7h
loBrnI+H5iIYwjd45eTsbZqN2Y1ePLunwLeht5D/SEJNrDvHeKM1/fJ3Aj1aFv2G
baAdtQyYzLMvGJn0hL3By/WIukAyAm1EraGsguICCDYBKDQMCaQJqbQc5uVt+pBL
xSqrj+6JQKCTewM3s7vH9lFPWjBOi63itJQtt+uhWoyWeWK8cHxeSb0mOj44qy5Z
qXXeBJNDMqQ1sjWEtNPkbsX/r1TbTK6mYbGsqgH47FVF4uQsJjzTCzv5Vi+9+iet
smS+fDuE3kCqqX3suY3x+hL/lAOOaN1scxVO8oU13437YkLNeP7hZ4VRcRgDI7pB
bAtLsAp3tSwtvqcUoJ629uCB7bKG/DHatC0P94xqHapCdz9vzZxsDqpqbXxFXMp/
+cWXqmIsUbMzv6i05C++1t1z+JRAgJTBk01FctvGL0fVfTHBONbJ0Z7Kk9jgB/Kn
jSm3OeQFAEq5ZPNjAMgForpOIi/AimZ2XtXkt8PW2XP8703Ug1h4MyTZKlAbbhBA
K4vfkhAcKSDdL9ZSHkqRF7C487cw1c9bc7e4bFiNcSDas/1AzV74Z13A/Uik7Cao
0w5+cDA46GPsZtYtWVpXmNYv9mQw0IE7fjR2XB5sXjwJaLLyYi0q8TmJrxGnL6co
syh2UAhC5pknqY76E0k2wCfLk0e24pQWTpFqAjAq3a3zl5NulDI3ambpMA5xVSXz
vZApNxm98q98UcoWhu7fhJP/Z3dEM75zUBAwqC/usgcN/TOA34YnahbcF9hN2WEo
4e+3UvehBEiRyAfJ/RRLDgESxbze6J9W4gbhlPMJR7wmA51N9MDZIF/qxZZ4ZiDS
LQwjR4bDcPM4XDnwOHaxYaFfTrSHfXwjp2aO+cerm5E42iea1js770LG/qxJAB1w
sUrV0GrcHQrTH+uPk3mXiwuppAzuY1rh0mhhZeH29cqJQPp3kJPx+brew89WIGzQ
IKG1UIhfTMlzig3p8uXsFEGygyAMRSHkjs+W5KT1jv7wZoew4ob3RvmRyoGWF5sz
siyQsnsyrMGSnMT8UnBiv0MBx+X6P0MqEcrOuWdktWx3R3x8GTYRpzW3oOk97GS/
tmLMNeILUMP90QOgvDhf20C8Z3R5aUOpKIMe9rt2L+8zpfkHduJpA2hlDSn4LRNX
WgocXSDzSy5IG21qkn99tPipczmH7cGOhApZGzX0ZAqBCyebHEI/g1VLUTHpCGjd
HdEsMcLDIDOvM5NAmc+TAeypLqeOOKP7cMX4J8DG6Mvn25RaOaqN5LWrZVU2vrl0
jUsxYEJ9S0NFln216BXEVWiNJ3Slroj2+wnf7uyv+AEyCmeuSaH7UJ4uSP6jjkd7
m8Dc5oz1Qle1HarsYA7KqADp02+V3fQGo/G+OiZBj59t6gC8heGwULL+LYOO+j1g
AJo/mc6vbfpl3CxsMpr9/G6VUWFITlfBsgG6ce8XizoeAurr2i+JpSXJ5c9+AciY
cVltXf0h70zB5tN54jk2yRhIYahkD8HWiydlrw++EdcAnno4OdFtaQB5gfVW4egm
dvu5Ar+x8/QsXp27FdQMj55dRUmSfA70LKRb7WQwRbpY+tUjhLImnKIXyGy1TR5S
+LCzb6FX/nBd+rik9X+uF0vbx2oRemRiubx/OHHVPrlAd7vHZyZRvHuiPHpSyq7F
J87KRuQN0g1thJCcuvGg+R63g7OkN5MllsxeVheAyyF28hSUxJnuogWhATH0gOCH
LKYqEcbQUW3keH0Z4ltrKpA8TSzbCm/58KbLxwkXLoH/kZBgwUcl7QWpm8RNs7Kh
pHlCVwuLPRHNhzj8wtPniVS/4mbFebnpnEt2NbiD0jsQBhFMyfAqf2Zn0MKiL7JL
Ibz8n+glJOoHuzVrW5zhv/vncBDhN05pDP+9sBeP2nTCuM4sjXlZHFyB4TsU+slN
t2vRNeYJjTZQCX4YvSg/vnVHl8FKv7cZy8C0brllIveNDHPU8TEdFk6G5oAMux/2
YOeJpfMrsoCn58CVcHMaAusov08NrSmrRJyO0nToO3LJbESuO+M2dgAC+LTE4zJ0
lotXsoMd6SjquHEdLf++GxUVXAzeOKcXMpjGz0am+5gUkW7I5u9jvf7YOZualWKL
2FuygHgf3fXx05GL/hI3qxXrcr+SwU+kaAT8yTEZ+DYXrbbm7jXOWI5ZexVGUrmo
QTA6Tvnf1SeKOvQsVM79Ae2bvhgYrB/iANKzcqB8Ihlidq4Cnin+FKqWB41R1Efe
T1mQdNkbuBfcRfVOBlLamq3sFROW00+uLWjB40Sd4wnhZm8V2TVUbHrHNFxWJshu
LzCT5Mb0e4akW96alzQkFrb5pqN2mnunW90dZIDeMGGO4WWIvAZ6k08v7Nru8lQ3
dza46bKrQwAIibfW0efmqVfajiuHWPHUYBAz7rpbq/9Zp6Jjn0HR/H8npGxH+kvC
Qw3PVqE6UuNxuje+HbUn8Qqgx0UextItFYYVMl2WKJFfBmDNc7djKAIx0b0RnLNt
ZBqS3UV0xfYTX9aSfCjsw0H/7f4tLikuhJYDCfz8ftxAAMgcQ4rJjZHunWGXhVH8
ldnMyg2AqW4P7zfBPNkdPW03HxEN4R77EhfYrwtOZ53u6s1jwiCe6tGack8fwZcx
nonUlr3M8Mu7fdZATL8ETkJkuC2S4yJ9Y+uV0zH32SNiF/kZ+XA8AvEFOVE+nnoZ
2LVQbKnmmD1lr7X7i3YD97RV7ixAK0i4y1NlaFEmZAF5VlfWkLq7N0m0DbMalw7O
HJpZfZgcjZopGnYtGD74UJLw3HsjwmmbPhsXS4kj6ZfvK504oEZEExxdQ6HdYpEg
XlpsMvbHHXKSZXO21k3mrngfP5xyYWaIrRz5vNlMQ6f6btU5VMBHJoJ6KRzsO01n
J3xvVmN9gbYWjspInlXFFgrZRaXXBellOKJB5yD6KZacSuQh9LGwc7DOaFMp89nR
R/UdVmXqc0eCF+Isq4MmOzdLQEt408we51RcImwKHRJTpeyuXKK8U9PvA62TePM4
zG599DDrkke9ul0Ye3a3DFRziw2MttVlEH3ULQLGpi1qYu+zIx4Y1WkJG6G2p89e
kkXBBkJB1J/YrjhO6liQrvTt16g1z15UiWLNIXWICH8FmUPkLHoiXtgGaraPIOm6
u9tqL30Pa6S1Yd18a95pcRt9hOZx1B8mdxvVEHelH4K3AUWAc04whGmlkurzY6Yw
oMQ8zsm/8drCL3QpskAcLBdbKiXl5EZ4HHZWKmZE/U79QQBw5R7qKWgnhOCP403D
uHmsZO+rfjNQJK6KAI2MGviU6FJ8sOTjefN7E1jyo3OMPq1jZqqA7PTxoMxi3PjW
amslMsLdpCe4bNP7eigOB0VDIflKuECmnnuL0uY+vn7HBfDsYHpi4r+0pl+beyvy
oGJ8a208eobXCGmjcmtEE07vpqyIGJ3ReGpGsS5sQ6zI+ZUJxpea0uFEcLmpK/N1
VdxVRKK45OTW/BE/MLxoPJt54XSRtEv9PmqUteTdIA8hju8kqqUhtgGk3/huU3ZA
w6pKmbdwaEm/ctA/4XhshCfVkNdWpvRxQVIlMY43zynh1aFOSuomhatUMW6kJ4Xu
9fK3Gad4CA6CQ+Mx0d+bRVln7y+8DuqWtFjwN/B9sONEcMi5KtoZciEN+A2fa9AZ
/lJc6ZQRQJbefTppvSFuY2INdpe2gqKK7NPArwfgGVU7n0FdaRZiSVisuHbLzAJo
01sVStc6bGcP2AxFlHPdl107//+FeFS/iS3WE3Qvg2bM3cLXcXSSlYVzZan7pjpR
dtyhLGc1B9L8PS9HnkKEZuRcgmLz/iBLaitSkxL4wwYn3eJzktmmT6oCX4fLrxT8
AqGIApYsfxBX8bywK8HKh79ZmAXaMkS7p/05kesOSWLQtbm/LAwFlBJkFKoYrz8h
A+wgXxG+7e+DNRvnoS+qZaTLvsRzxwncvJ7BUxlu51zhGGITkRuHaECd4XFC406V
0HQ0mpqkquUtzKlvK+STuDx57OKSxbu7LNfnJYUGIjSC+kQXIpThvP439VzrG2gF
SSir59hTv+x6Pm2dQCTyqTueU9zrkBhmpj3uMpP9fy7uMGIBEEqvrMsjpsKRHeNP
rjBVCBTx8yNum1BsZesL+VozYYffget9AvSH17r6dNh0K0yKsNa7IELq9DETLkA3
o5hyKue3RwfyyxJLNtMyqWNQ7EdEKBVgQK7fRceF6Ckp8YD0U6xkCUW07N0hc2gA
E+tLHGq7hjY+3el9DBNZOg9e/mIyrw96DJ6fYIqP/aam5L6vTuvQCLA+dZGphgI4
qXV/lyYer2j1Wtdww95uWmXrcvPxjXKhYarYG0QTPxb9Nyq1hOrNqeSez2PJkalV
XdxyAHVyvDpZ5p2UL61HnwtIU5nuAMTAAQg+ND1SgDC4EC4+UwhgbXpCvAdSoQVj
scK5YK94T70fpi3fPyXT2Autlko8T07as1fX9euyAvzQgQLOd1wExGSHUcwAXZWf
1f9nRCckRKvxXfj62WpZ9goqh3SmsTFhoCjAxWIC8CeAQNexb3Q6PGopsS0uqtrq
y1RhmEkOPDXemS+dO1gaLh92bchIZmXOigv127mDuj/J6wNTxPgS7hFemop/HHsW
v2J4aQtnqQ5onH1HKm6ntqFYP4KyON9tSr5MXPzNnwq7g7Fv4s3Xmha11f9XX6vz
0YR17wo+2a55oBEBhYDh0gSaHWvFLpRqY0zgfkQMQXpA/pI/pwtoazKIoncmB+h8
gJ2tgo/scsatD0QEPsEUAPTjMhVWSHvgdc+nvtwqtzMPjnG7FxmYjaGkbkXCps0w
af6Gm1826cte1SFsx8pVHaUfPWbVHCinVRKGlMw5SgFWg7Kc6iEHKaMSJ12MCgZv
4B7BndhmIx3sU0lTUjHxtzTDooEjx5GIzuKUhWU2gbxmEoasQTGBUMkv7rUKgp1m
00Qh2IlOCu0KrIJI51Pu6Sp0ZtDxU8O37rLORaYnKwtSh1GYeIVEIygTZ205L8q5
vltRnkC3JO6M2Zx6dkYkWmH8ATyWgQ3bA5yAKN4MRdMJ1q5BD7rW39cr6y8dWLE9
SqRvg3N6NuyFAcRA0+fpX/+i1DLi1db36DP8Plt1yYK64LHO0Y+WpCFtlKj192ox
0Pazsbsz+Kda9nQ1uY4aHcKDtD69VgB7NskGcRMqriNZhRmRJgO2/6rIw134wQrX
D02bPooWWVJNTZH4T5VxWc4FXLjGiqEyUy4wg4v3DOls/NP5gYLxSlHzIKOL/B14
L7FRjJwGAkeNUa9SUYJRF4rsbx2jdzuMLudf7lXGOWxOKoV01tEtRHqmRybJDDSa
y3VJfweIuccU6l9EX3gBGZJWF5QbXCc1VnK24ACX+wbe43+9kqm3HADeSH7GBeao
NsPmhq/djS98Fqn6EYBBV8ybnxcz5RtfHs5h1irCY/uBql+Ay4DDbpPlOat0aHBS
vIyb96Wx6E7/XOBxaCA/RKfuszHa5UfCVLBTknk9a9ifBnmINLFnrpSc7IcO9sX5
0GIGt28TVkqeGYoYnn+NVExugCs9QSrYdnriB3vj3MRUw6RLCT1AGmqZtUU9JeVZ
uWkC5/nvoMXa82N2sQ69xyK48O8gndOCJgqE4k1bpCLb/uO1LFJfqu8onmVs/UrD
T4cgCkxdv8f1XnKqSZBlX9wCprxMSQrNxjF20g6mPqz5ku2f8GbQYTNZqAIl5vna
OV+xQTcFCMigurv6L8S3GQiT6i5bx9uK5rh02jk7gm2LhTKEyukCCev4wDtFDvkG
cD3Fkc59XPJFTOPJArPEdz2kVZHduSfTbcyR0yXvO9xwD3WI8ttOoGO1Wq5Ru8ck
fJrOdjntqpvmyMC95Rd4bgjJKxCL5sxNGvQ2vhu8QYM0ZDSqEHjTjoXTlSVZEAm5
cJEcihxNG+mUHWeJ+RvF1usyY4Eppwu+muTvEqXcL7yLnt4eR4Prn+SSVoMlvjWv
C0QBtqxC3fQHKXqUFpx+zWIUEHJxtJ0sVP1K6wis9bPaf8pVi5gGoG2OoJHKi2V2
jzl+oQpoa9Wi2Vn5oJV7RHq1iIDVyb6M0e3yZ/tiQi4aVXsyfhzwvZRRE0DBE6e8
pHtm/Dae7cpfYS7chWh1XtZ4x+bnzoNDkhgtxlnivd4GvxrX++v5SQsb93uru8Kf
eTEt1XOqEC4PU11tuDfIUZa7oSpRNMUhaT5u0z1792iIIdUW6ngigfzi02b1r0hC
P9nrew132eqSTq6rD30yFaiSf1jFoOLhsx8qYL8ueQOb1k/7mKsOW3xJ22tRwX4l
AaqX1xZDDtlDcmrmsisB26zhDP70DA5hLx6U2oioRXJiDllJmNp5IrNqCFixErtl
Reu1hvfdugoaD9Zev/mpcIS+7PiBKCUH5fIL6tgyOttPd4Ym3tfNtIKB3PB85mIw
KgUpih+MWBsKpC53DEBsr6Ot/m4up6yoMUJlv+b9vwdQW4iWzNuMXwyffo2SawTu
bb6FoHLcufdj6pymHysu88sVCobkKUPrfT9sBdMYthCogNMmUIw+LFZH2akn+mws
8gqKbAi0gXylOoIzjf+2QwGAEsJ2tqqklbAlfGC2F7Jg/jRzexfqQ0TkOplt9Avz
2ILNtZU+LrBBnIYAB1Fi+Pxys7hzUBGPvpkLMqygRVs2CAANvDk1J+UFpaOxhhwG
g3DqK62wPlct5cRkAnHlCP7wu6yQvxatnC4JldZbFQ8buObDWLFGbxx+nDyj2KaC
0GM+Kvtzd2vUs8buDf0Tqo+31LR5qPdmUFl8SQD+ErKGyx8aAv3zP2r828XjKGFA
IFjdA9QWLAcaVHVOVS2q/laUiLFcibMztTx6+byOOtILDFrUwVvK0LtJBTJ2xNnu
AWuxMbmxA9IYIjH/k08Nour+KOs1fmfvVu8UgAesQOOasyV2LT4DGvzO2j3fWRT0
RoPJuaPsdoGZMr81oVKnhJ9u3ZSsGjfRDdocz0xNHAEAMGXgMoHO+dAqVFW0v9IP
Tzx+81GfzCkMepE7ZzAWNG1oiDbbXRXs+W64DQSmnBPO0QGwtjITJYJbdF/dkpo2
7j2FcKwAB/S2dvg51GN8QU+pm3iLT6zRSnEsykTt1J5N/6OZ1kJwi0iOaR4bQMn8
HDja9hohR8iMg4k7C7n6DhXU0bvu9KaVGvLDHp4tsiOzpIBv9vVwMiCacUdBCquL
Tg7FqNhMNJ7ib6nCVduhyinfMe4XgL2wLBJWZ5fUwbXSKkjeVVh6G5unqXTK+4zq
WH2UbWPIHXSxvTJFtUJL4LK5L539Ij8L8NUrrGgxAIVGevVCXfJVbgrwMw9DHOo6
QeZR36SkzWp2vroSYGWqqb6LINROrbG62Oj7XF2Ut6T55Y48aTkDfsqTl6szFGvW
z2e3Fyt9FLSmxtazBK+9DfJIMe0+JwinDCxNvHmbTHAOgaIxIs8KC1sFRBCpCT6x
/x7TCRdNVp4porgDLTaCkBNua6GRc+FAAJRNVjqJgEnA0zCmYvFpGmSkJTfRIfiQ
LOajGhoaMX4tKP52zehZDzuQo0ewXX2G/DKsYqFM6PEyF1v/Vn+Hbux6WcHtQ1wi
5EmQ7EDc0a4DYPr0heYrNYsPkjDJ/cvVHYLvk0ldP1NB/9aEM4X35rnIt6uAtFbO
sDYJ/PXtRFiFEz9/VEIWywfdrEaCmxbepCbvK/jvV8GFDV8pCjjCgmZqEeCoKY9I
jW81G75M7toTb4i76MsZsLUuDbj1iE62RiaDUSZacAn8q7dkXaf65MoKAzFQtnTd
RR2vVe5POsoFjFwwcLvY7bCMAhKFgEtgZCvzp6ycjG429zHDs2YpvjP9KfKytnlo
MfmDXYSexyiRgZ+Nnkx3mQtr1+0OltDHNqi45EcPi/r3okxnR3MDfqBu35YLh5UF
yqgNi6cOQGNZPgNvLENQwh2zOFc5a2P869JArh/vBOfXgUaq72tdAx1isig+R4hx
e6AadyP9LcvYIKeYzXF9e2uSUPOjcBaDZeGJLB7siSjjb9xpuEVCQxZ587NJFryC
5yRRc7nVQ4VoA6r7v3a0+dPMqOJjGhMnweishduEXA9cWBiCYHUj5XbW7YyR5GuG
2UFOuQPo/8uXp+xwVduCgSCy42MalLRWZyNU/QGf02IkOVf1ndQknLnYKo0t8EJn
JK0bL4n3/89Bk6sfKrr5Xb4DI3Te/01mtU0JH40sMEsaKe/KE5iNm1gP9w3mdKmS
HbfnCrcVwZoDEYhP6YLKOGqL9iz3UvFSPm37JLJyqTpd1rCGSL0tYDTOeI4XkW7U
NfSqle5ESfPV4bmz/r/xaxTPNcuztKqYOZLjq5QpzeQBmW+QOy2I0X5W1WuLNnve
BArR4uojI/+qlNGnO9yFAKnvqVxQ6NeNNZOckPljK4qG87xqhMxCzfYj1V/+nxM1
hjRyZRUQHxC1n6nehasnUXoucIUNq6kvMdpl42nhNhbGGqPr+9jHajsA39ogwHX3
f5q94qqx/YQ8n5Mw40/tsxaYUsp2+GjwE1N264rz8UdIFQkF0PeJOImy6J0icMjF
uXoVFgpe2nwpv2BgylxrM8o0a1nosYzYSN2uecz7YBx98xRJnzmyj2mRiEkrfUDK
MR1gIT/BHbRdS0zPW9XVMmzybm0NniKLIYI/mKwsTJOGYk4P/3JCqhmcsL33HtQb
8EkSkzSuk//uIw2D30xSYFak6LH2MBtQrjNmMcztvWLnvCIKiNvMAYXc+SGXAW+5
9xCQLROHLjwD8TQmx6jHjlYN8ZyEn1qdz+XsXHz9TT/NYSV8yc/PVaNGhrXiX0dI
yQfOvu9pCD3eO/xyHToUcwCIh58lgpdya15hTLPUJ7r0Ro7B3cjY1QkRgS7m1Etz
BDLnQIndNxNzyvUKikiZ0DiabUZnn8JXnZl6YSm87f8AnF0jsdXkUxCd8O1ZjWhC
Y4G1VFdfhVvCqWJhD6B17Yoe6DAXU+pXlqtCMmHffGWvPA2E2lzyp+UiJE8NGhrv
HB0hl/uSD9o+25eoklDQtANkmY/MiRWJWDY/jDmmzVYYduUE1eQ8Z+6+WF4sYQYp
KzPh7wyXWrRL4hFaRtQ75pOHnk6zAW/i+UIoUVJULwxeV+7DPzdtsGyUErNJzSPE
TSqHp3+eFfQRCnuhwf4uJVEOsFg5gJPRUijApiGQykMCxzruEnlVEcD8b9SYNftO
JywVY71f8Z/kT9TeAY8cFZzkIXF5TjJ+52zlK2dl7aVHoyKdbMfpWOc9i7qySFiw
V9/mytQukZtBzd5Y83+kijdZMXVFNGwPhB+OCHQJI/8W/sIB3kaeM8AhEM9R5D6R
bL5PsHGVzx80UxAwI3ALY7Fna5A7WzT2HWYdXQoJ+2wAANoCWh9CRyJrgz3PaxIg
9ZNH+Nd+1cM6gYF2mFwyBoaYkguIbt6sHl8ngGgo8mSNCwE3XfNL48HxVgi451fm
I21Vw8yfzq3jQts0WPbZLItdB2lkKOQvY3TzePG4xiWZeMFhZrbwry1PRUGs0s8j
7uotNLuFzJfAVkUy1sRAFp2wxvfEnGqZv5q+Dwg57l9cNLqW46494qIozgT1rqcF
eIpHbuq6PrIbETEZwh0lSi+yKaKSYdjKffb1pNmYfk//s+jyFdTNXt8Apf1DFC95
fmA1soubbhejDye/CtWgeMt2PFT0oCyWGFN3R/SQXDpOxIQ8BvuLyaEEUXux7JNg
F1DzZWsVyYqJELeuwDeGhZEdulChqQ7q4Nq3JHloHnYw6j+7RcOEkMUSNu/48lHD
FqhbbyQXN6xq8wnvfJn9C93bfzHSQFg6WP9JFtCPo7Vfi6AaA8UweMOLZav7/fK1
JqeGy5tKfAqcL/RK1olofkZ4EE/rQS9NS2Zb4yUHrNhLWIoxOV2zKF5IKlQ0H1KI
3Uw4KBUdLRE08w7A/o+16v0oaSPel6FPl8sFc5CD/auD2ByjCvQp2Jy1KgoCjU1A
ahZ988A148g59JtuF94DmQ0WdskZqPCVnLjgVQIXTqZLOUQ1t/OV4C+LJdZ+QtIl
p4sM6WihyJUdY7KAZuQB6YjNdAnEM8fVbuGK8zG3lYY6k+5vawqFK8WuDEuUfNyl
HAu6xN74bB5QAib7Lr8OqmhYms3mrDc5DvMMQqMdyN+SVXecYTZxeZqg009RULz0
Tf3YC2YgevNH0P/rMLQjatfA6Dj8xjfDitphtPzuah/GTPmvBK7L1Nxgnz366IHX
afV/VykyCFLwU9/oMmpLXsdfiEzXIEIJBJBtu5Zwrgj7FWOwVbLbBP1K6rcg8yXd
46zxnFYjXNZkvbjsh0vHxgDlUdkLdv4gxidDAf3kFnpWQUmMZplNnD5IGLYeTCpQ
6c5nFMbFVdBVaOryXMg62ZPMyJYXbgpPs9LcPp/zpyly5iTTasA4elar6o/dO4S0
v3sTTYHdxHI7Envqxc09aAV5FQ1wFqSWhbTCfe6i4VBepHYq0RwCTtElF5C1bUIQ
q3f1Xyzix7Tzt5DLq2Y0Yx54EiPLAxCWj+YyFuDcY+W+yf+RZkc26yoZRxQD13he
uxt9sIpmZAzNv9QYS0xUBC/aEbQc6Q2VdReu85Ge59BElfxnR9lgrCXvrxB+Djab
GabMh/DNWI1+Ivy5tj+L8Cz2R3xhwpzUjFGtrWl/NpY2fReRnE/Jw3pdroIZVeHt
tARbt/b8ohvzpLrKUXpsFha/gJSuT8FbtD1cBB55AyWAYHTKwidPmPxnbVyCrj9Q
0Ssls3/2dRTiZKgJY+gMKB1B1s/tFRF3ZedWpOyosu/JX5Xc+g1mqQ9heT3WtEvm
I2Xa8u/kErYlXeopcT1DoWu5MrLfQ8NQjmv5XoM9xl5Nc5WvqyxKR+6+NpO2k3JP
wA577HI/G/xautjozTSGT03Bpj6XtTlWLFH1G0x2nNkxFIhJQojJ0BIv5PrOjI4Y
wENb8Ae0+hIWMSvQwAucxKlXd5l+ZVuVy3Iij2dHzsFY9OlLfZpG6g+M2wi/FUs1
5u9pysBNQ0B/xguKjOoe+PXxRcaz1IVc+LT0f/l+LwWMUfb8dBgjmL75thXWRhNN
0X2/SugrTPXtYgusYU5WKnTPV9l8LSnEDienbiEp9au5wOTuShjhfAZL5W2CssYJ
aM5GMe6cSRQybyNpmomCmKGbb6j9M4I9tUrguARxeD0hnhNWBSzAKJDEETl9yZeI
ipZugZFWJJDR8hNG0ZmANxCrXBJtF/7MIbskCS2fVqvnHj5aYhxmMbld73PJiGEZ
Cy/wzEwNyCxpv+Bgk95pX8kvac5AKByOLP2iPH16cBOC+hI1VEOJWkG9H76eOqGh
T5XftQhctqHwwUC5rs5XjoDlHSj+OefKQOQqW/qAmTD4YvUoRPx1xCzf9UEkUjNb
kBhyI+zfgzgT7LKnPWfDg9P7RSu2DjqzZXqqUeLfX4B1XvitRlOUeeIvXTlVOIcS
XtlZsUPsigtEVoueRjMbISGPigTnaNlsQByj9UPFcPyuE5AIyC/NtclI7iEpPOM6
8q5eXLWqcWGtzD/zIW3QjmHz2M918LLIAJI3gkQPDICU+0QNy5fpfoATyIfWxeyD
BW0qiZxS93YVhvAMzAZ0v5eoyJTefdH6MAyN9w6cOKPO3smzJjL8Cfkx8fm8Pcqn
oCIPABeZsmJwmM4v5Oqs2C7wZ1ydWTitHJFD5FivJBe1LMfcyTyoziylbZMx2ceE
vnHDEGbgOPqcYv2ArSpiGekvI0qx68AhAkLnSwLH0ZEfOb+JBkZGV7NR/+H7fO0m
vy8F22wklbOmAVN7ofP3xcFzNPydwvRmpWUFSy7HRzSw92zqhDJk5T1LLm1a+Ps8
TnLJ/FIQAfCIIOU9GOwoIqRoIqaxpaIRC1GO17F/DGuTwlLmp/8VaDgBGnVEWoQJ
UKnwiaPNDCfSRtw0mEvXRcensdPwIkDJvBtUDU0+IzSQDisTZYh68+9NEUvL+oot
FdnVuBgXevByxrkZlXtMFwDeyHyY4atHxM2pDpuLa+TtAzhwVcPCCaje8Lq/jJl5
uYeQ4cHZaJU7ql8oZ203xqTPnUCcdzM481zz9oSVhXkM4nCQSYRUIqyqS8IvMUWA
qkvMhoDFZlYixWgcx+h0QETwLBP5ayMID8K5Z5dLC2ena2IgHnIvvopLQI02qVTs
+no/5rou51FvtIa1yguOgG+iKoC/tSdWqLCTeK+xOzUfCO+E7b8I1w1uPAD6XuAA
3wKgcf3c9H1KyL9RIO7qcAh6foSAjNcv1bOhnMbM1daV0VXsOfeUvFNsmKdtJcK2
OjIM6b2oXGS7eHox5McZj/dMk+LihgDYPlbQs0YRqavE08zvbJ/jVy9Ta7eFPW7X
e0fCbFM8DtaDhBPxVM3IDOZlIpsXP36HZRHdwWWR8XKJRvSFXNPII/EcNMM9Y30F
3I9JFItug7stS5uMhQTmv1sVyls3L0IySSIpGEcUjqhzeK7aC4T3Ii1tLfsbY0ks
SPOpQ9vgaHviHa7B+soTIxYU5kF87FkUs73Gszon1w3dFy8LH4uZOVZ7BcQ6pvn/
rwyXhXkW4Vmkl0Gvs7la4L7rZTJKYPZe7Q4eD9orJZhLlg7Hbq5FuL90KjTmFRi9
r9zVpaN/80GkT5FR4/i0tpJonG8j1TdcvGn2IhGmWJdADvSJQRtcjOuYhsKwe55A
F4RIc4FAIh3o+VOT8UEIXTzVZ2MTPhONqZ7OeHIF9Kjr42AgbwAmRj03o8paIg84
DtVMFG9NA3BrMjQvrHNkyCGxTlJj9HF6WP/8Tw6t/q3QH640up59H1NehsGT9dqj
CKM2ezpK4CTruVJ0j+hwnwvpZOf8RQIX83yrba3yu8zfX1vNtKNUx8e2C3lkrCC6
DDcqP4ilMyNiaNDqihlGXlhuJGGAJ5OZAccLSNc2/QpaFXZhSuaKEtAydA1QN8LE
txU0baMR96foN94T7f+ouKtX5VRiqChI+UpDG80+hL5HAl76ti/aJ49hgSGqAVsT
7TQjbHHNhZR5OCdwaNKbs5kz/x/AE0xc7OgpTUZRKjTWVYw9QV49fsPvstCdJO1D
Vz4sVye3kdUdcm41j1mPdzyJVLeOM9nXKOVsskEKf2hTlx8ywkHO5UGJT+puMTBP
sJFm4qqXS17SdPQ4xsnLZ645UZZloZN6qx7BCBBQH3SnGvalCzwsMPhpTJIIs6Mk
xwbnfh2O+ALqIkLLpHhug8hw7K8iKIn/W7RDXA47eTn1bb71BMgrzrQ2ECt1GQMo
p8nkKJLxeE5SIBVxkoo9LNN07ujA4xwM/loVCgorc8aE1k4FxKB7FhekwXlA7uKZ
oGbpJgqtEX3xE7F/spMIkU40bcl6D4GSaTi0mYo5VWe1UJxdeyVuwIDDjZQHmGvQ
f9NYjz6flkrvksdwEDLUUFVQQb1ZSwrA2Nsb/jGK9J2qy2EVz50tXllJCSnhrR9R
4kWJOWTWI0YlnyQ35GBR9vp26/KaODunl5zx/cE6a3nr2LCA8CB/jsR9bws+11Qj
6/JR9tc7vNPqISrguWyv3fCTrBexBopVXQZIiFr2vrHwJ/EGZwvRBbhoHUcxRT0b
wn8jBK5HlxEjUz5PVHe7yEA5xW//8S9ZRixTWTv72x1cOTp4L7LTkKJWUJAS7xnu
vQXxq7iUPT0P8tEWLqwnnB33/91c+yG8cWrmjRLAEVe+i/6S9JOt3E80BgkdMdFO
DIJ1LO0hWCVvsGQ8UrFr8mAhDBEkyEJDvZ6I0nEVwxkL/YTS2/V6vgjYdvE+K2in
JkkK7Qc33RMa+v7Xohe4O6ZACZd4UvskrvDQFI1PpAWyF2OdWrC5gJ0Z0cLra1pT
AOb6D2438/H3Hj95etfOjAQznqC+iHJcjYwH6cwkXp0teXa+VZ1mcujQGIENKd4o
bgPs0QKvMKNzxMhLuvCY27qiVD5Y8v5E4utWbTwpXNYiO8fHH6P1u0uedIj5FNtk
hxezgu14SE07vf/klLvn+ZX003WlRhwEZfic8EArlMw1bzm4ou4Ks+egPi3DyMf4
JtCfFKCRVA+yZzjR9RPFCXCPX5GrNm8IyupDIutjCGVrFReNk38J5BMNKWzULhqq
q36HFBW7ac622C4XS2SrltOVOeHyT72Hle1GblRsCcG3R/5AXt9jlHZQl8wVf9Wp
RmtHlyCyzRdzvvpAT3fi40xR8m7f0dBdGKWRIbRiUpbXuxV9ZKziF+LiQjU1jSt1
CCBDWaD4Lwv47/t3gWK9RkjGyVmxs3sBb4CdoKAutlRsvFRa6D5U4puHFPMQXsFS
83ii0T9L4bZjza+s7j+ofEqo/axNXeOiyqvZbh5pmxhOvBCHsL7yyZN862W8XWy/
fltgxfENuSywAMzRpfo0gVucsMhO7+ZtlvfWP8upt21nmSge8cQn9cmXWxMm11hb
RIzheDcFeFA397NK6CJ4DDEK80u2PxTq3ezgir2H4mrPHKO3/5Dl6ML4OVXNcFmm
0ZcQ2AwVDByiwNbNv36uRkfYPP4sbZbNv0KKZqwenvtLO7WFX9QhNSBM2tfqYeEj
qQckCNtWAuUDrsnBaOeb0AUNcquGgb7MkzwO/ihUeOzQbBpYw0YhSksmc4EEjo8H
j8kN2uQZYyUB/y/XhJBwUy7JzPm6IXsqY/w3+8/FB0Df1By8FyL40iiflrPjGJy8
XupON7xUbRoylyY0vlx2W5Jc7HIWubfEKxKhZCA+MApLSU+CnBjtGl5GcKvLwh9C
btm1R3ogVRGB0xMbOKK2JWzaHxc05y95qrS1OQobNyxzahPaN0wTVvKk4Zc3384P
0ybXIw2RGUaPwKGWApLQGAO1G254BtnKUL+IcN5m7QcWW8g3T9NRA4ld5K3+DFPA
7Ll7FQNVywxRfslzRA7YEDQlPJZnjBj4nR6IfyJOTvVFGhcHJgdYwFl+yw8yWAFS
cm7AEH/J+Awo6QF9IkuoQAUYI2ZIakERIuy035+Oz+1A+ndhiRN7KTDlZDVcfNn2
v35zQf1iPxpVrYOhN2S3sZKRLoXSJz36NWJ1fZe9svNTdxkuuiU1hv0QNI/Lp7xU
7E2+WLP9b8SGYeV+91vlj9XNutEYb8qc5O/jPjnGUrhFsZXLDD2uGy1EQ2GxHBYH
7meMJq96Fv8ZSjFPLpAErfEdfX4zktjEJCWZ3jaaw1dh1J9UBu3cByDnsTe2OVu1
1BRkFp4NZceYilwxC56WUHA24L4QIe6AhmFLWOWeR1MghIer14zN9cL0PXnTv1NI
1a5vmI1eDEczoD5Ajci2W7L2Qdh4RI7A7Eyy8ccRvihmUTtLzrD0JCwVLCQkOtwo
f2D8RTmmFib8FCNXhP3YIccj4OQ/ZtdF0iGiSIZ3QoAGbDHJFcQu3FbhhUnsEAxY
w3CQHbFpKrvVab2QEn2oRWi9rSrnB1GcXEg+N4L+0CgwnemhP+jowZtJ9JxQe4la
zUSsLf9wQ3lo9timewnW2qgv037+VytMJOdBPGa8BV/xrzGhjV9o4dWMa12Tlc6S
/fURql8xbrB+g8AhQvOD7a2qQCMrW3hTOfibMqiRJ3yk5lGnQ4OQrFYDF6F/HXAm
C9vETwI1I/5yv9AHw5a4SJTB90t/vHVMYLUO66QOUoTU/ilvlpI8edi5pZFgS+8D
RGRvOKukt9BNKfSVBanTdq2oZJvK2Vfd2q+V7tlGYhAX0Ut8DWdxSRVgaV05++wa
1VsL8CNIPd6b3y3+GkyF0fS5H0MHDmeKehR4x509vmSeQVO9YpJS8o9K1SNgOQ2N
qHnm8REN6tSLqYXlPaG0G3sPG6GIpRLBt8xttfTn2+9Cx8d/EXDIVpmZJQ+8fp6W
+/lU+hFxBX8zLVLcFbPBFdXvFpS/FD52Y9fb9bbOh2/F1tsn8jstr29FpFqjbJ7X
or163T4C7o0K0CnCgl6DWaKWPYkin0HNcOji2NSSmXATalK5yjMj/GLJ6FL6EjdX
vsDa0QjNfEa/7sAaAhGcIuPFp+Pfof6G8i3QGm85m1EJ3UajZrbpnXqG8OQ2MY2e
zSdI5nCkM12WhIveV5C0rqMi8B9Ym6oCdvm7F1AS+WdDcLpvhHtWXxMjC9l27mKj
/GJSSUl93RxozhrhwBk7OYSF3fOmm/YR38YUHLZvo3YyANNgm+H0QqQ4HBdvuyHW
6qinRFxQAFwxSuqKGm6QM9jRTj7Fk/EInxFTzrv2bH1WRG/zboTzJ8NI9GaFfXYk
dmHYaHQvFW8WkLDYMM9xdEc7L0nsi4T9PVvJoUoACdBadUA/L24YNcsGTkUO4noe
pUTGQnN8Borbg87/En6E7/tKcfEX53xJEJsrPgZtk2Ty2Yi5K6T2q1UsRglTRqdF
jwtTVFedlhLuEqzndYgCDZu8SNvIGxi9xuMTYyoGhb36qoZSzMCK08gcN09HRkdF
y2Po7BCyNM2IRVw6fT9slu1nT65MBJAQXfvZogDydH8fJtHzXJd0kqmY3Jdg/XFh
BgriK5HeI6xvnOFO19XmkobbvdQupAFaNAH/Nx5Cjw0Nr7vkqE3fe1wiFoy9tEGq
0QnPsA8/NZEVm1z+7WnfgEMaAIqCShNAwTnBTHt/Pfwx2rjyGecy4vyusE2yrz5u
o6BELBegiQ/p8Kxmp7cvVIdTDs9NnL1lu00Uqma4QZ3ZhK3UUnlBEZaUuxlkNAd/
jokaoIpzgnC6eBlw6K7O2pO3Lc3bkIEAzHL0H/afi6ZHN3dsr4HA1ccxo8yKaO9d
R4ZWomLWGLhSyqDkMbbeped0Vm6s+ctyhg6zXzSL2VuCvJhwBGZStpsLTP37j0C5
6f2opGRvrDORROn4HG+CbKoAsgP0krUc1P/gmjtQqNCWY9enbekiFqryKWlCiRIj
tHctIBwo6PybbyUyhf/4NMKStnLkJoiOAbgftZ5TP5+xBUPa1IcLuKCdTkbGEbn7
CWPlmNR+YuaPceAdiCC1ECB13abybVQ7Im3icDx7e9AvfK4rR+3TlhkUiNbgYjUn
Eopo5s/PTpb0q8CfZayylpE0Te7rYjVkoQOGx6dkme+Nx0IfbIVzx5EGm6/VDqtL
NuizUzfVjPAPCx1aYQ/y//aM9hOdsEXHpEPNlewckjmd38QYjTIPeOZvYpo6jPPy
BmYTaH8X3HLZjbumCFF2v0ZyUdtCn7d4muBjEPViaJrQWCG32osaudBtQek/UnTL
RJkNeE39aozjSfp+L7vkAJ3DlQlGeCPKGQ8gq+gkyqei7uLtPR/gU2C8mEIZI3kY
d4vsa4YHlzRUgv4bzmmXjQcToXdjqTyohI0s5IL3MRKTEhuEufD/qX31n/xY+Dtt
Maqb6/gATh3FyrXaDZ76w2KdnXkAJTs0suv9U9kpK4DUaQ/ya7ajPNtV98dJ6pLJ
bPK7HXrbvfdaywNWJIx3PEJ2vwi3NnCdGPpanINrxgddb6qH4cvN2YPLVkcKbeod
ZhR2iKEPJHdbnt9HpS/a3j1TEGX3MSs4xPUO24ombN5aYkWetXrQPBtVkArhUavg
KeJvFz1PRRalrhk9AlHMFEY+WzSIIehxn30MHQz/mjDIvbfHlBSuvwMnxtblCnzW
qmUGFgSi4I8CF+fg53Qi6NjfFHxvMh2zCozmaWEJyCHYbCjMbk6/bGBo/GL9SsvU
QmitwVA3RtxJ7V/LsQYH8yYlcwtXxxr+N1dGiCB3kcMkpoCHKyXOjxF0Nwe/MYor
Q90L6A8f7NsjGSKWPCy64ADhZELMm/VCMYMI4+I5/nBHgo62bSPAWBJRfWUTATl6
RwhmKRINfBk6T+NL71MErJOrVXwGSFAUhtDuIIK1Dhsuxw4qM8CZUniPgzyFqkPz
Kh05NqugWdY1EdFGJxtxjtP4rqipOE4BzB5kyDUdsBurAlDAX7NUL91cVQCCsdtu
sDkhAeszBsibPimiOHgU1lRMdW6vgPdx+VltdlafcaW6HJx6bOvzz428WkConisZ
vzTFtptb1bjAJNfyavxW8tBvSmkDeUPw+Ew4TsV0SgqJw2+cOrLvupH56LaFlvyi
V4wMDkQlwbO9oYKHBRGHvhWEKZvyoHs1SgA1XV5Nb4i1Eb8QLqx7VAl+s2g2wlLh
PbWr4W/yGfpLscwpXHAoUQJuzS5UpFo4Czf2TupzCiD3l21nRs5SbEZ48fp7p0MK
yfRan4icfrIIq6ZFFvjUtWOLQCgEPmhYYYARYDcNZUOjzW9qqf5iAC4yWvzCudGg
hY1sa4Pl4Zmyg457wlbZOk4e+pQZjYVfvq3qIO+pMlfAVlNn6t/lKe+J/+n82XBj
RZTfKNT0Ko3NxQg39YCWngOV0gjzZxR+ympik/PbHKR3280I6O6i7CTA8aKkltne
xsdPj+mcpmath07FmHevOqEy+qVBvl2kUy1w2dmWM1Lt8Cy46+UlzROxGnee5RL2
1e0SkOwpcshq8JL84OGqoVMhTcDnCLjfqwULeZcOLZioWAzYtZ5KC/IZBUkgt4NF
pahfRquBfdSBulPn/R08ph3C9z/fhmLwNl3IQOjlFiyimbQ/cVEfDgpflUhbwHPS
NcgDOUTzuTFEgUQYNO/n0TJTjI8baWvr7eW4odFeSRRNwpaO7HWWqgoSaD6MuU5b
SVx5vGyUY9r7mHQf+gmJWQEghHdLMQ+xVuzP8OWM837A+lfsCyLeQFj1LnXKy36G
Dp/5dKOlt4yrU6t8HA6ynoCHwbiqV8TRnHyfaXl+f2qWCEHdx1hmP2K4kh/gd1+j
7XW12LrWvW29XjlWxJTv6Wx1rip4KDHHzTHx1/GFwmyP4hbqvFptAHmiy5dyysXz
2JbeiwNlESWk4D/QBPDMPHaaN4REwSIClklhqT6zEXVY4GI+lk93eLHEy1MDrIY/
p99Uvk0OdPRs7/mi/HoFzYrDrZUFYMhPypmtTVQbGrmRozKH/uaLkYn/NTXKg8RN
y91vzBX3x4unhKH1xKdm8hiusK/rRNjQIx67YDOSZlWCvijNIEMIEMD3s1ZlL+XP
JBBchuv/TYYgEKkbXa6BsNaVld0l2+i6m9xivfu1G2mzkvTTDl4kcciH/knoouj+
WLZFDSHsWxiuM0YfcwPtvAtup+1rM5B0l3ZmVj3oU/RxIKok2tinH0Cgpuf0dz/T
y8MJNWHLnfdv3eseoE3qEB8Kc2ZX42rrMPC/mUxsUup2IvWQAbgv6hOJku8sXYYO
F1aN5RzO+fRtPBvwYubaFQxwCgWWynnkGB8GXRyJq1/KgnpOyX7CL8r3dSN1xq8z
2pdC3RSyeGQ/nWwO3UNJNnNu1D51qxDbexdhkI5W9CSDSOnjb67x1soeM5NRBBfo
/LYrMqwdd08HQOF4n6rZB7S/6ch+lhVreZ0wuLtLJEehftsjEhbd21lmr7DvHVzo
ywUfjWpjv2rRl9ahdJ0VmvcsZir07A02JTC/eR0h6zvnQNwiX0mNAHKo81lfLcz8
0d8La0Olc5EtEg9RRE/Q1NprPZDzgfcElUVidZ+CnVi8y9KlzlxvNdArzyv9bkbL
PH0xzW4Cnsk5kAg3oMgU9w1Jnnwjn5NDuU9eJ7tCuViZHvIJZJd7/3j1qoXZNjJd
ciKa2HtXcma8ZCLVP8sS5H1cO71RES9ElbS3lgtZuU0/3ccvAexiJJLKqkxQwUCj
HWKA8QVVouFgIUHoB30ljkPPCPRafbgMEe3bY8V9Qc1C9rc6uWz73IHYyO4vTsM3
vJ7nvwHVJEwhEOPk9xDfrPLY80rGvPrdxadcO0i1INF/bCUrbfyF+y0egZPVfoub
WXzcPyuNgBWzDYjCykb1zmC2pBPJOSruxd1xJXj4KEZH2KpBFsSN9TO828IVhbQQ
R05X7lSqO9UGwB4Q6qa0ahz87wDW1Vr4vpRNfzzOmXDVNyJrp8sXyqG9K+rUy5H5
6USPre9+WxziQ0hJ4k18guQVoW+0+j6PG/c8J3GjqbsrQ/5484lpl8nNWmfK3voQ
5TBIyARUpmodapIPklguBK317SO+7T5QJDT3Ki7OJ5k+a7Kv0IltEjh6gJ+uMQIR
YVJoPZqq/oB5qumQDu2Bd0+xIAR2lH1zBUEXjmbV9prty6BSwiUPrp5xE0XCZA6k
i4ZlIJPRlY0vyc1peD8woHZ7+pWfK54f2kCT5YuU9b15mR9xHKf3UA9ktO4pwOOH
E3iAT3jCR5ENt17D/tf7F/gwcB3bpk6wqi/6N3nUIYXWnkQkC6nme01TLSKxDA8G
D6hnhG8AUyETQQoZ1uDhEVBoCHmwRon4eBXE6+AeOd20KhPvlrMDqW9ORTJEYYxT
R0r25gbXW1Eq8Wkavz2MbtMXkVotSJZLnPzTI69cCZziN+GlBWZEtunwJmnXWFr2
FiPuNF33McRV1Q9KNdCVC5xeyAJ2CChNnKgIv6w0Uqn8OVPVO+gAEIAZD5w5dv4U
xnvul3Pv7c2Zy4auIkjrLDeOTymVRuzg3VCEf0rgAzts/idK5NlctqymAsO/4Yoj
sXM/gD0sy1IglYmZZE3Tmr/AfDuyWMaoXfj6vjY85R5eVmIEYXL1mqUS1Gj9CswX
d10v5LN7qM0qhDvHV2IhZ3qZfMKndtEibUIKgvNPbQjYW6STK/D3/9XX/7Ey6SC3
79ecTxluecfeVnD93jqaoH/IhA1z5gVZEMWg6DIIs7Ib8i5D0Z9Ga8kHxUGkLgeX
6LVrXvyPfJAX+ta0okC9vsZORpXsXY2FJZmxkiXkKzw9IhYl2qSSF/VT89qct+Bn
qQnQplZFQVLF8huOCTTF0DsNQvEHBygkR4rO/M6/+4c+j55t97fnWUd/Pj8ZG1A3
gjZ78PSgO0QZTL6O7BTaknsNIDk0fUdo+wNxq9dkfEGufEV64JAi8+P+4zqKAxlN
i3ZgqP8RQVIZkFAZjMRteG4eCGFMJTKGCqHS+N9STtrxgWj5CkfCS3O4WIC3OtqV
QsyjfWvlpR10urf8G7PFY0CD6sSry72DdBM4qAh3mFNlMYFjbmFuFccoekfh6Nsp
ureT4p3SaDScq6DN2lM7pKjWjQ/zV/aWHzHl6sggUvIB0ZrBa74meobd4NPzkeAc
maO/AMMn9C33xuMYJ7XFkT+nTNwmiYVMvx5U+a7K+JN6q0m54iapacNz56vWxIMn
DbJq89ViCZeW6xSF0jnjZY6F414WpG9r2GZBMNGIxjdgGQMoBz5k+WqvCXQ/RglV
zQzleQbQGLzRz9JhOcfg/T5LlmSQdDSs7odqxZehT33YBLschzaFNurpjXi8NnaD
LEIe8wx0JgGlRtl3YpuB59rYNERidMx4MJNZTpvQlicKCEXXeR9Yl34FOpsz4PW8
rPN4jF13iqEgyVj4iCxRCbeAKSxjF69sMpWOJ0rSuc25GRlMHi2Fd4Fc/H5t0UbE
3aJoJPrB8wACZyBT8gXGvao0frmw2xFgiJyeiVkeDZircmtrzQt8sUpdwww05vry
jQmScfznrQmfZH4LCOzaZJfUMoWDMez7NYj8LAEc5vE2Q95eBPFl87Z5YqNBY4nd
ck3rqbxcE0nK5fMyKPf5tZgKTPe5DHRXnph+QCgpStSQhdUITC0oI04IMPp6DLr4
c8E2iAoRdVVSdOg7f9nfOTQh9yvX4ynjFZVF7TW0gbJLego8HfC8XhcVsIxpPA0O
u/MevLEea4e2yBxeFuUZHuanybbhKRdYnY0zxpMbg+iq9Kc/gHBqJnYe+S3jtyNI
75my/kZ3Me4HXP3m/3L2zKmLk7B5X2XKFPtrykJ1rwQjT+ysuh2Gdx1ZETpUFnxd
gqwYe+0LwVYCBEClnVnnOPr5FBO3zZedWCN9CV7KPPe489VAEaTclLFvAKPwH1cc
yHTW3jct75ici1K4Qmy+ulcGHGV+mGf5zSA0vuNPvguldf1rZe+84M11DDX+vWzR
a8naRjNqyktAGJzyBGbFV0Cp2XjmU6PUos6mSQFQvcCYv+cL/chdLpTlW7E5upmG
zy/tb6JcCyWDpFhZJf06KxzKM+CaV8ipKWj5NRe4ce/BkG0tDeOw3q2yMecF0T15
MxRarzS57WTPYCWq/Y1nsrSRY1IhasF71rvwazd0ysgRfbKZ+mOKx6yQO+UGNOFE
AYFnXWv9jX1RXr6/iONt45fLIE8VY6Z8jtm/YTKampF7O5DKlrRh+J8fKJeAHKOX
zuPDALIVy9bhSIG+/86q+FnbodqM9F0QEZU1OsPf1qhllvLq8bKMthy/IXm++drE
FCJQzqD4HZWEIhcENmMR+mL/7zHj1cdc67RdZLsZamNM+p+t2ywwtQgmQVttufuh
PFOsd8nBB7aeVG4hD//lCMcKpkMJPVduDtDGULtlsbA9MJ8RODPJDlZuf0Up0AVb
GOBpTlXLWHO5MdW8hb0uf+h+5uZUuYSIS4AjMg3y4CCfllJ1nTktCuIkxnBgth1f
FflGK2MNExUdO7oyyiLZjokAwQWFlWNa+46G6MKCCiCqB6SQqzAsZ5TASNHRBOhP
VmZmgPggrnrx/+j33I1V5XqcplFlduMtfIyp0argATGuixfVICONVMvZxMqNoaPF
gCqBxopCs9ux+YcQ5KBJJu0BnDN1TDWZqgjvxmdrCkOz94cLw/wBgBfD6AK3SObm
ZVRR3AfXmRkdSHDCHDqo6z1F4ypxf1aE+OWUx0+cP1GUn6sr7MkIIdrgZhlz9EvY
N/DHMaLd6MqwhrDtEwatHbMQI08qw1QUvzj1TWxUa9PAfl5SP+Z08a7hTCRpG1l9
IV1PCX7ty4HkxrEcrK5k/b4zze2LJi4D2ulAYlxokYVDUiJOqYLJ6w98QgiRMd6C
UzUWYc8ohI7g/W4Uz3Fh0q3Myvyi+l4y1/w6mPNPXQ0zwG4ujLcktmx6vcH4ZDDY
cEDQyQh8Zfm3Bs4vlZRFL0JUQY7DofYzxQ+AZuDv7ifLkzij/VVCqxjrOXQf+83I
QD02TV37TzfB2hdQ5FwbIW2V1Nv0XmOCKzrweSAi/856xSnMCtYjxxf1H74yOJKT
O3qIaxulshDJzMkuaJR2MtBJhf1JgUCdD2Vp2xLS+seBw/GuGK4RWioM6xs+RRZu
Suz8tBkvPqfHFheW2qhLZRJS/VBXW2o90/NmYnMoWKV5b+7WYWtrYARO+JCGlFy7
KO8ZiW8ZwVJYJm4QWN9JK1VHhkbUmJxqmtY3xxlX9pcsfBfpS12o0ApK6T3/biga
t1rQBbSFg+wACFCM/kn58EI1rEfSPWyxC+6ldFMHHBS7FWKpC/37LLZ8EOvkyy+H
EptazsenTSynJKow+CIEe5zwyrLLam4+Ja07D7Jb9+sB1aOuAHeg9sDCjkqkXS5q
6faZlUhKOW52xsnhsjD/E9cqmqy1CQ3bJzq1tNq05WxTFfcXw6c/Pu7q2cjkFhD8
cB7H8bHm6nHMIhzDdWxDkmETc32EyZLp6N2m6KDdfoHgFSem1vQwJK4AvGSzQDer
XWiCLPqzVEvUPe0mPsKL1pMBaJbnoIsJx3/HU1v5VCOCBFD5a9NoxVzVuIttE13J
wOV9QxnF9XcXwW4XzkYTQgiHnu6odzmnfp65aUxYYVtl8eH8AdbCM5fNPJzO1MML
4sPnUI9y+UZCJEvefqvQiKRnLOeihTKvKWEcAbNa6fVOnFnJy3stGwrrzytakkYN
j9HyxKlmvznzjyM936c/GqUF19snC9x4GaCaIePFxrATGQ/8T24V0cvEtERbeznv
FtAGwtL4UI3YGVjc62ohe7bzeYYH5i4gyQBS9PVUJIKgBZtnsECuGGb35wyWlaCD
67S3E8DIrgyoGfxbzv6BUgTse4oOhtnaGOvVWPWDiEO1KA1b3JwSwu7Y+YzlN2aN
sdxKFp7vV9Psns3A8g9boNrTrawLWFzK/18eVUOfVJzggZnTEE7xCRZoZW9Gd/LF
JlEtuCApL6rwEX6NpD0VrRlHhx1hczrT+ozwrHbIiR3aXMXQIlGqzuHDIv6Fh8jM
5U1+fkWVTcMpYZ+AExZOfpAOvq48XfDRi0UD1eYn96JJErTB6bd3fmzh5LRkFtij
BJiY90sA9aoiQodSIR5mbxQWJzLQHrc+B4po+XwAr36jNFptbcU8bQHR9pDo61qF
j1LkO15lCQdPggLJc0i2mdfwvrhHIIw8SQi7mMRmszHOpA2um4iv9jleutu3rFTs
dDlUTuR0jN9P+B4Hc7T8irTAcAm0dILQwp+8PnsOa+RLkn5yYuBE/fHJ3+pT5QJ3
Vt7V6THF1OF4Z2vI+fao+YZByb6WVPSy2hewdeyAQJSgkoFhpJ6Zzd5B+n52uyTl
Of0YzDt0Mr6QvAI91UCX5YMrKQp07yeo6r0vjysRDMEH+qse06GxBZiIhxsaoSpm
UGpVTU37w+/ZsFxsj9hFnnkuXFZavLMN/ZGIO8+SELKVcZupEz9COqY5hWpvRG6w
ZE7zGZqD/CkK8vZbo5LcgABnUDBF+vfjMijULyothaZF2faEMzfiPWRtdHfVjqm8
MAZuQsxo6XLCUwdq4YJqkENqpFgGBoHAsEwKf2Zhk9jEfELj+gFugxRU3vN19EUY
vLpHztgStRcLJUES01aM9nNNONRtT9gA+TvM9oH8Zm6+CNQ1LPk7CFIou8rvsV9n
5+NnxyjNXN1gPPjAfU730z1bS/8K9PJHAix859N3GDzikb4g7DC7MnWcpH/an9Gz
gctT+x60o7GrnM4syk2NSI0BQRVun88xXpw5wRnEVa3/zWowjEpVyR+0zPvpKSIe
MiNTjAU2wzuB5TSdYwLmpctt0BaIJQsMxslacEJofP5ViBl/u7MkW8Pma5Hg1Neb
jiATz5c2zIkag8wEFh5mKBqrSMmUhGynYmntEAm7jHl1BEoI9uQ3oIIsnd5K6nqD
Wny5AL+u7UzQd7ZnvNfBggIY+qHYS02BKGBUDiOcT9WsHuDLSp0CsGDxoVmDu99R
Htp+sy53p+l9GudXfxldWW1bb4DbLn7Va7KeOxHoPq8/K9h7QBcAFjml9biF52WZ
LjzeQu1zTP5JbRHU0XrZob/rK1X6Qoa5lzZzHl4ihaNMCp7rvKD/cstQLUYlOy/m
J/m3JT6lLLLBM+fYnkCJ7SbSJGGxJCLZo7PulJtM3hYRJVC5qBo36+GjDelIuxFs
g6aEqpFTSGLO3Y2Sd54Xali9kSiiZbTDsELGvXlPYYYQyGtyHv+V08VKo1AueDg5
kVm8dUh6q6IO1au6qEDLe1xtFt+gjoGKle4W7CNm7lxtfmVEZZahfVF7KNBvGH+n
WVa+xLqlId778cVvQdcSl+YSI6Icq/ytRAoiEW8649zrgnw3Ywlud87dtQ+DYO6D
Nn4bCdsLG4jCxLtLTDE5MBT5X6UH3HCfUICREhzeyFoG4oiAafyMTJlGmq8Bu7qg
R3dStvTd5QelgHDVB5Ci5ojnNBxNjUIA17bf463JDrg7vIIJ3TMV2aDBf5mDgQ51
p157/rlGA0+61Jq03Ady0LFNfpRC6Q2ZB6IaHVV5WeOvQwcuDCVm1dXI734aojrM
wi15Ezj/659t/3iH0n4ypT9WuSKtviqCsWcbzDG6XLy8FKoCK4cmcgNnS5idYFLw
RMXJnGl0z0MzeqG9SQsy2LEkn714ceZpjmb98ZUIjjLofV8KpigAQcNLKUoiKH0i
P1BnSP/c00k7AlVkR5A8tl6R/xi76Pzi8SrCcTCYB0DGIbWkxPvITF1N3MBpn1SA
ARXaxcfXf3T3l+yJnF+wNX2vRh0qkm7XAbQxyaeWiBbTCQMSgJAMwOMzbfZGJS0J
a2glZ0ONHDTkpyDsRSDveXdKEbAcBvagbwIgXeL0Wfx4GNcClXnJwdDvw1Hw7SOX
FAnxkuDPbq+uFDUZ0sFkFepFBdi/WbE493bEiH7DnBdm7tOdl5MOnkbcfUCTEzG6
+WtoWyus7NpzgDv4QSbqVPgl7pah3TZQ2k+k+TSNIaBfhboRhIIB0G/uwGmVCM4/
ScTpNKBezkYf6CvV2xQDx8y1LP8m1A0ONjR/IoIablOhrmIp+uDT4U/lRaJs9v23
QM6tMRK2JaWfbv3bYP/hE7TW0kb56+DmyEDy/KlK8JCW4JesDfjZeIEaZNZA7hPi
U6qLcGURjyP89MagP/XBI1HDFxhI5B3H2ri8/492PnH8mRr0TEC5u/y5EIFbjNDx
bM0CooAVhn1GbSWkwfNP73acacNA938l8e2uP24mV0OOVNnTlbXs6jFTL80xt2bA
czQJ8MBuaUc8t+IJj7+xXsqDQPoUaLg3DejgkqTM+gXMNDOc15kW479nulCy/MwC
/D0fhG+1oP/4lSQc+5Yn9CLZeqyZIR8YqahwlftVE+EkmlriEqSlJe2tUwxa617n
1LVjuzQRGydnQANreGIRsBITjUaFV/2qqGgOV+Wp5FWAukDK2An2eRDd7o/xop8v
42YAc05im4I4CKnLeLaU3R1yxu/WIfEzFBI61WDhxZ3VVDHuzxVNZ9PiieqQ+bVL
rQv90Ger1GStXUSJWgqtwtrVfK2K1nwkepfBUUKkY37eaG3HbdQ727H782YqJUix
fFqPEyOmvg3M/SQoT1scVvoGEitpSaFfz3/+RGz1aSALKI1Uq/EzxGjM+qaJhSfQ
ol33EuUufqZrRRZ2SqZVgfmbFNICBPubRyehygsXgo3aBMRy7i6Q6czlqAha/cOd
LowYVPdzURSg2c6Zj63l3lHoCwL3kbHw1QzYKhNQSLhcKgxqYYMz1uo2z8tCRnw/
/2Lv0lT953P+ys/hQkl7H6/M2afdbSmwn4uPrjCwJvcNuit1R6+Z/lEVjpogYONw
hc35Vj7DIpTd3Sn4Z5usLQy9eef2YRHhb2CIjpJMouwUXL9Dqg7pH11BTGsvBv52
enMDY9Wp7XjwzizWyTYqU1rRSWyukI8rWUzQZSV39YHdSgxhotqu2Jmqi0aCd83a
Ajyj3ni7lWgeRQc2/Va5uQ1/Ov6RdHO4txK3qTrLpBIhXPoT1g5GtMcuT9oIo4zg
sEPOTB99Prn+r7irJ/dKCGJ+dbM7Jw01KYLRWm45XuZD0B/4P9qM+OjQgxer6Nkh
wG+dWwzz32T/C4fTU7oy+eUbvUn6yMggB2dEJjYEQ9eNPiHEzNpYAFMQ3hHyhSum
mElw5m/gK6uCHGc+7/+VIuArJXOeM8tm0f14U2MRRZGQ+b61ZjG55Oddj7MLruLl
p7dbS6yi5BZmedNQKKgMGCGIHt37oTyNgLtvLTZQzMnBICRSrighp1QSXnb56dGU
j1CB/JMX1X/m+swkxGuP6oLx1DkcSF7qgniSQIwM3mxRUBlnl2TdLpTr2xU12++r
bdb3OHq/o+7nbZ49VTSWXWbDpcuSgUIwtfiH0k/rli6HnlKqA73DKOM6VNuaYVwV
fNazvJhA3UPCG2zfFvwrxYf5BevQfCQapitCZKj9hFF5GwzO0Hqb4ZQuq80gN3x0
57ntr6+GiwQZIZDaHgrLSZynusEvundo39wYoTq9mo4c194MjYiLGu34eZN2pqje
w3iRq1iL82+yKUTbd9G+spx4Ik8rE1kyhOxfghBW8DJVOpGWouPXLt3CEO+u5rh4
5kzEtuqBnv2r7xCSYn6/AT3sd6kuq8lovX8vsChrA42WMU3HCEU6U+Ejx6LWLDwe
0tP3mIyWUobqpHTse+VPvwnsOJ1ZwW0R5IUh5lto/0jEzfsrIL9IH9Rcpp2dbHYP
fRaY2DRx8KxeCIdfzs6BaSa+ODJxJOPmYB+PLsc3RUbs0YDUIjeoRgvt0U6Avkkf
tItT3VMNiqrkC9Xt+gPfTWJylWLTgId7aHqzVr9yZ8a5as87G7lK7+IaGxJyaEw4
LN4chVamNFCrNB0+0GVjk2nhRhg+L8oQ+tac3MCJhqa3tlsUmI/cAmzjdAzXB5D5
cKF3l+Q3HPLmnsnc1/IS2Jhsm3dg/Rp7E8AKgmbQZxnGX1OPpKqLz2EM9yYmNlvJ
qG/R/q/MZ9/kzsyXd7MkM4xjPxlya5XwP2ldSCId0vowXA3KW/5GEzk0lVg8eNUQ
OuFGfj1YxTGq5wV107BWgbioqwSGnPi3dZxZpvU8bdfNXhUz242BUZRQvRVwifL1
Yngu9TXYU+qea+7hJsGjoPPUiOYv3ZuIxrDc4xML7Ucep2HpUshVYvAp99lBEoUh
N5TegFt4fhOn+arZ+wwwMEDcoBuq1s0v231FV1NIKBmz/EeKL1xmViTtX75EfRtk
ZKBYZGR7Frb9lRSedQ6pIkauoLt2Ch8EuHHgyIkB8SwFsaHZ3JtYTNlgfYJYYU7+
wzcZLR5HhzplFER6Huaz0+ib1Bz6rcu6y8zDgNlbO62uX2gq9VIUyMHLeIuzZDrR
Ho8Ffw0NsNGtwB0HZ3rKKga6oNZqJIe9tw5OhgOKuW9FbCuDF1jSHGn8yKrJRruM
7wagY5i2qaukqZ4r6DtIb308naOuItxRBP8LZp1x3A+K4R8+9RskPirBZnZOP/ak
+cKzsujIUtOad8qf6wafCjiO0n0Mn6zJzNRMWKmMzPq71hQr0sugqjqJ7Tqgtvt0
C36EiPx+6pCtTzvxPzRT604cPko/5rQvU/T48I9cyK1inaxn2G5fwz6BlqurQeDN
FFcyhi3mLsILfvP9LBF6sM153YZODjY0GGAE7SsCrKRKd8jbsxbwPj6JMp7Ajd3a
k60Uqbj3agtYnAbZ7yc8NPFN0PyaaNTd+W73zOLB7OXP3nu+HftL18oPfU6X8leY
MUzH6OiHNClOAahknPnzkh2hCGexaZgMzmnQIOe5uDHufdMna9uvpoMk24lRFH1+
AACnjuGE6q742XJ4UlvSuIp/04zLTBimVHWVzJTfCvBrj9XQeaXvmwDsJs3BQGXa
5/i6WaEmv2JIwNfv3aIFZbqfi7gSf93pEMOrsPRqiDwBncIfJeiHPDgDNbvuXhR4
1RstyQUnAEVdI5xneiINgQ125GYJtAORxXSQhvLit8TUpAi/HUhUy78AEW57SsZg
Vw/jHVk3+tDIeDHWCMUhKM0/cpPS5RhM658AHaDYdwV6QELC8Hu4SWKeHgLQFFAd
lA2qI6DHIOy7hmZLEz6LpUS6JGKty4BeoMtPsy4NI21cakSP+XYT+xAz2afaGpuo
ufupkQxtHvAfFtT5jfgTBjVKEg3Bw8MVxHArbVQ/15a14Jvb4Z/YjUzsdLEkd8/3
WRG38GgyK8LcY3Tby8tXGup5K53EEmIGFDcB5+pOG7tjU+qQzRBGEmfYzlVjrCYB
mCvI9+waGX8gIdVMeINsbFZT1Zy369YgdQMXkeFLLEmAh0o/B4K6iLA7oqwHOCiv
HTTGxSBWNObc4JC5dcxJXlu9naOQd4Eg8Kq0RAOQCiryxJS8hneUNiSpVkTfA1g9
/aDPFRPqlImpCZ6LTU5q+v6MS5cYuSVM+VIAR/+i7Oq34F5XHrueTvV61uY4mOtg
I5AI/JfgNReI52pHW0u3UwGfo9+h4Zmj+seJCDxmxR2LSolsByn2YxmKeww/ONh3
SRPTaJGvvW69NDZ98ij/un+SOSc6o2Vh+kA6cKysav747utfuR18qR8sCQnW2Yos
5I7KfVzEZNmLTJYge1my3EPi69nlr+sn4uuRR2iH4QxAoQhWUNj6kazJtF2TycJs
S/noFPj5P6anV2KIb0dRcU22mrkuXC5pwlRDbohzCTcqd9UatRoIrIv4t5wFzOWv
3akqcn5dcQDBaCvSvPMJpW0rLIFObPjft1wyacErlmQopsDF7fkJ4tu7f9Uxbc7n
YTk8bmog2xMSoZbqwlm/JTVT8JpQWtd5je3FqA3tlQ+sNQXUTGMkg8YHxCeMPDmO
oOykYA0XxnFZZFUcuCze2GqrEpJhEUzDnc4h5hDeUxdbTjCctKaYlK/Wbsdmlmy5
fr6mTguvTiAQzUU8BtVdsbg8ixfOYoiwwkV9daC3o6Gx3artRdIh32QFm1YLAwui
vyEU2CyCvyGe9+j0aL58KiZTp4K+qlZ7DgtGqOleWk27hFmacrzpAgNlAp84hnS6
3ZhtcFfwLzsTFrgn5mD+kSIziWHbZ0I9dqpdVgDqgmrw/elCehkpRE6dMOROLDLr
IGr/TGhaoGTzoZ1I4ChQCQGFfpbDw+WvQ3OGxIkAfp69z4z5DE5aAGgFmYAQLXeP
7YA5uM2eBmB8iyX3zVEovZMqMWu/b10adxtJDfD8pCf5Qzc2C9zDJODAGEm7SQlj
bxm72zcH/Kzk4MpAH8PwbILdOgY/Uy9RfJoGnqbybgmZM6+CMfVb6pit/OESJOp8
VSI+juS9Eq5b88PeGqjRy/Ok1bnT8w0yuHJ8c3XD9jPTESmMcUrxkTZfuywH+sZN
2zSKCBLeuAnmE7RZwst3rsHaIgzPsDgVQSluqS7cC4SmAIvuZXgeJNPfki2tOYV4
UhA8n3ebtn/ZP1DPnRIT0bCbM0/GRYF7aQOHMKsJ26HQQi7PQeExI/MOLc3T+nB0
I0E4rQSnuj20PFiKgW64RxPlJCSIDGjcjbQ5zOWZlyATpEasZIPnL3XX9T9gL7h4
R6KyZy/qLzLxk6HFi/U9swakL6bgaYwo+KDvqLe/bp+0EY7CeaarTp9LTD6IeN8Z
YgWCrC40u/gFxd9nETfIkDFnmvG+LOWkMBkj4ffmmrD/N+rsRdqU5BjUomKW+ae0
AC1DVcvTrPnxM3KoPLK5op9ObpMZD26m4JB35SPoBuEugrSUmcKoTcfNVBc40JSn
4XQs6HR2iSpvULU97T0ToZK64DkSTAXUd02hArScm++sIJjdiizgK1vHZ62ATRAH
YQ1yh8VuAqvtgHOP1wmys0GiLLrALFXk+hUE4iWok+B/Yrw7899HxFo3QGxZhivT
g26/52q7+F+IOGDnmFmo2TAnxSYuRNL1SOEB7s2ZbcPpjejUavwiYioNdq6dZufX
+yayRDGmREUXzBo0dCuO+B/jlgm5udMFfd3KFfD4esrZ3yR/8x0ooTfFsR1bhVy2
oIcLw7Eslhn7LSBy6FAgW3NFIO4RHnrYJq4pO7TfxkhdA1C/XBUlVwecynFJARL3
Z8KGgTj196Loe9LncOQ9h0K4E/kbD+Xt17fneKKhs/a9Buid0Bq+0+bRdYsWJjpG
w09N9dqjIM1qNzipN4Jsj+fYqhhCOilzjydqD+2yaTQaHlV0pFKRqi2cuL0OYRq6
4H7yHFMfUh39xgqjRKUZRGtlIqSLibGAIMtOIs52giIklU+F86ubdVDE6pW0kvP7
Bi80upLEcRpoYH17t1WkxvmGx6MAXZAf5oiCPoXksi+B+84tlgZTzrlO9yfRuaqW
7RUAY+XbAAjgUjpDjfXjqdAcJif4DrGpyKJW7d1LARDNolDmbCAutC0NC7YFyQDe
CCQwRxzIngnqnOnLy5XiQm8VCjUiJIaPP8wEhrx27w7UHZtnO2RGfSTLnthO1C30
6lwg4WzqRPg/WsfUuVAELkqbQrwGojpb0RdfHoMQnOP2+H5B1IbaKbOoVRA7gkBd
nljV9g1XVv4MyxADhHohYkoP5qcVL5MWWp45AcSiGX0NpwtVT6FfMSBRR1UZ6jp/
10uOyC51B/AlB5uNVr9SZQWH2BZ+KrJFQ9rNeUDvUuWyEFo1V7RvS28V7XhoitCt
YtJeH8fGNjdbdRu4GO4bk+gbyHV3UEkmtDrf9f+PnayhLezmmVXBxWgOwd2hGSZ7
bU0Xb0790R/r1GryRAIX9Hc5OdevOkEiFaRlWhAlX6UwsgvF/3mLjE56PAm0xDpa
NlfNdzghm2WIHVaHIFGBKySGyagdvd1CSnUTs9UEPL6jbj2FLJhee4uLddeQy9DB
AySi4/5pW3WbwCX14I9Zwe48e2+nrmW9b2IWznBy/anaxIlssBjuj0n9aO8ts3W4
DGH7uBfneQo4peAs+nzjO+6Rrfb3dCQFghPkl9MIMSzu2iGV1UU9/e1edFDNY/CQ
OJbtZcU3vE/Bpx8XeiIf3r5QE5MQGSafSHCnfF9DCWldN4W8dGG5LZjQ0r9eR/8Z
VXfuQLv658p9gMC9wfR2poehwxYNBw1y80AsU7+dwONO7UG3IBZuGbVVe2IMaZGI
jy4k9xuE0Pm4wECvOsmz3SohcGPquX2BMtZLJ8dK/lsPRqFSOKDBViACVLh7nqKm
KC+s0P4mGaXzz5cGOjPO8NpzvAwxzivYY5ZZypdkk10O85sIMHzLrG9HsXqKCcnC
FuB9CL8G9MqgKDFb1SbZkllMRtuEmwj6Hx0PITYLQ2oLWhVj/3ba08Hp+uLSS21i
MP8ujtgyaITePwaGsEzlPCRewSZZXK3K/6NijN6cF0DDddAnjruNqDWJ1Ief2/Ca
Cgar/meW73SCRESQDzFCYBiQIPhUGs7Z2hsI/ji4pYV1bU7Cw/W1dRp4n109Mfyh
FfllRDfsIkMA5z0QOsCBWR2Etv0xuv56HhoCkK05f/miPjhvXoJbPW2FdIHQ0YLa
4/emPs0xnSZGX5ib7eUdkEQed581aXOcrJzYqPZ2fxOM5xaUKnLNIJJkMrLjvOn7
Pt2641V/jOgZ/7fwJ5UDU9sMdFnMr/c0f+ymQgZFnIoXGBUEvnNjmz5TyAniXRCD
jUr6bFGv2Yuc/44IaNq8LC3HDd5ovoSupNxulZKYj6pOTTh1QjRPWSof7YMVceg9
bdaaD/FddkmtrEs439MVCC48ZOmA2bOA6vX5uO3Cq7i/ZiFOrqyHxQGigjUJXtx6
kpYTigFqM5SK4PHV93pN8uZsQdgfu8pq1V47uYA0SSW1Hc323NIZroaaTe5GFaAE
OCfTpYoQi9gtmq87tiG84A==
//pragma protect end_data_block
//pragma protect digest_block
RMsD5wwSAQdRDwJe2jPeGoZ1UZ0=
//pragma protect end_digest_block
//pragma protect end_protected
