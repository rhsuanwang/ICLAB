//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Oj78Y9V8QO10Wa4jMOfqSLO+WOgFNqYtxzyIJU48xQ8HSajH5sIll2F1Hv5R/UKj
4lufzlQvJf4zoEHR8kECIvlmrJPfyQRuqXgK02wrZP1DDFFxB/pewNS/5nNhnB4d
MHjetd1rzSkWMqrDw6VmNSukwmxEzsJBh2DKlnCw2X577vF7Kxc4NA==
//pragma protect end_key_block
//pragma protect digest_block
9+sjCnuYI+aJYUJuVE1PG+50Om4=
//pragma protect end_digest_block
//pragma protect data_block
f9gVRg+pxUGUrdoED9cDkBINGaBe0BF2Hfy2/Rhl54kpIGujK0Em2RSlnblzizSY
A7c9AZbVf0fY802THsAHA5BNTIk8dHThovLyCDNYOt7jjMiWj6NWIhkUAVukEDm4
OG490R75an3A9JkVen003o+H/kJJ87foNdvKDhO736Dgn3lvi8N5yx8+uNS8ZZqO
J19Bdb6jMEZIaRwTIz4dIRpFpXF+C+HUBKB1EbHOBPx9ePZV+/oGdAxJZImV/jpA
rmj8zqMWdIayCJjtQkD3Ed8HsVkNtGtyHXeX/FQcqh3MKgIgqYKW8nMWRfPMiB1N
Tx+l4r8+OrE7YRfae5gWWw==
//pragma protect end_data_block
//pragma protect digest_block
mMazESElb73aewpFwPJhSK6jG18=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/E0MEAbVt/4sm+ply3wV6uI7xcC493M9pLVDrTK8wWKBjZEIKSJSDywvrJfwiVtO
OGNFKQFEwBpfz7vGf/ENWpXOuDDNzECepRaTCny0opFHtsBn2F8+KJHS3XjhTswr
W3FjhxW4jZUxT5uq2URrCwJpGLvlFtIi2d2v45Q/WJRc0NlBSHd2qQ==
//pragma protect end_key_block
//pragma protect digest_block
c7GCA0M1oAOCh8Y75r80tkh7Iw8=
//pragma protect end_digest_block
//pragma protect data_block
74waes0T9TAisVfRdEZY/nwwW5q2OPrwUb+ghx4G6kcG3qcW3uusfhKO2vRprjxf
t3Cc9RPpjHfWuH/kSlVrEJY6CxCFjkd3xeN14Vy2UcvfDJjn0M7gdcX43HKe3gD/
E38cfy6gCaBSGEXDsyiKbY5YqRjs81OJEmlLlygE0IbLjiutsw6izVTF/juK2K+k
hSDvJbXcv8Rr9rnvXjumJ2BlB29wIhM22Xu2p9Fw+dtbm0rCWgWmWmk5AAHY3wp6
Rad0MGXxAyP1OrFTXKnh8CB6S2Z5hsxIhnhen5mGzZJTL+NEyqbQZDsUNqBhOHjp
imYHeCWssp0tiijq7fo0Bg==
//pragma protect end_data_block
//pragma protect digest_block
qcSAPYOmTkGo3SqQ0nnKxn/MGNQ=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
p4/166h4nNjLDcW6UawjpWoXm8coHrxwRSO0hG97ku8gtpf6rdPzPHdi59+R5p2M
mg2whOfGyZ1LzeRKpf0F5Os6Vinmwy/H9esA3d1ioWeI5OSCnCe/k/yj+uNfKK/B
e+n6znNmQmULwTItbKGw/PV0f6sn+hmYmMBjkqUgGsmv1Gn4VUkyQQ==
//pragma protect end_key_block
//pragma protect digest_block
kbPRTKhafw6efZBpT+f2vtveqpQ=
//pragma protect end_digest_block
//pragma protect data_block
FHr3F9kGvNhpXt0DsMTipVM980eARat85wxBSAuaVAsvCigm9JVI5g2NyWOA1uNh
N0jVHJdQ6QoRIedc9yqqFiBpAAXPSt8ksIIdLnLZsXdGZ+wSjiNYaMX2yXZJ3Edn
wEIof6FZUABTLqFAoKjFu3F1Mv5puRXvRVprTBqsZta8qgpqi33i8kM74UxHOE+I
swebtLAOmgZZGW1x9rlUTa3unFs7HYQuRfQSf0PY4ncSuuqUEwS2kppDArmXradJ
C7WztWKDE1CXuYLJMa77AH/zXAzjUE9U9xlszI3eVyWcB4rYlID8tGJxdjwEmZO4
jDQN++Blj7K4GJwIrW1uT4klTEnsieLMocBQERocAI2tlluG3TD7Ni3KVQ3lFRNr
3OGrAE4VP7PZvR1a6m8pUHcruP1Zw4zyaIQJzIrYoPuuxIBdXmffx0PFeObLGCJg
O/hYTGA7IkazU3nb+l7z3rPL47b1z3mRlARnOOAFsw/n1vQ6b55P81jzvRp/2+f7
TTCQtwYJCQ2SNz7syTEE449FGvpKM8tTTiz7qgR26qz/un5QUSuMTXs/hJP+LEH9
WpCr6KNcH5HUIIs3tvHdgweKA/fL8ryKGZbvCrKS5KE3XFN0999JXDpbO8iygOVc
j/EB7sOvz9+iDicdGV4SMNbg1Kk8biWg3Zq/couqlW2NbKBhaTVfRMhegsAqympm
xcXxBeTQ2Qo1E0YirhS8HzI41GFVQEcK+LpHV0U92TX4a6n5ua/0X7LXowPVUdGg
gEnfvfxzXeN4aTIA/LHnw4zMg8IlJnRiYh+sWwJUP2PbGF6XNMMK9b0fgvZETktv
71UHt73Hty88X0RPKe7Q6nZiP4UC6WedC5QfM2a1m4awEOotREGUGjjS4YLkU4GY
wnE1jWfhzpp3khdBeCoYSwj6Y2SHfiT5MW9FUPuewVgbr1Z1p0A971rw62VQFIqg
+8NCHK0cg7O+AxumlnuMRcRm5QEBhu7qwNMsf0m5opMNzjF8vrPCwe1Uff72STAT
OpI1lJc4WvNJw1LS0oWkDlEAmJIX9axbQYfXNYJI2MhJu38zZuAcNtf9Uh5QFUZW
E+gCzTMZ7jzY7D713uhsCvv82UPXqdBKNKQ3YeCg/s3zTn+Y6UBaSV3WtcHmu+q7
yt0hMbIfle7VP0WiUL+Oy22qpzRwDwv81tcx9vn8mAwMOIrpMH7xQ5c+1NLUJYwK
nQ5dwd8HBkcuT4Tkyz/ocMCsf6JR7zXPZr0rjtpCSqmNZktFbUHBcqVwUnAL8scw
Hgmrh/GX3oaaBjFhkq0HedlwGcBUNLLvCtdUFpvp5j2PE1FhhPLDVOHfgOCn871i
Y6vfhnlayGmkmGP/TR426cvRkTD7VEHA8Y7FXR3MvvsjU99PuUuAoUUFFBpoaRb6
JXA9xZxgM2z3gRKsI0rWTUh36VcS0PKn6MZpoT9cuOo/tkS3P0mNcvFSStPhFnfb
lNeg2kcUpLdcF3LqI6gwju/ISUfJIp1PESKmmZ+f+FnriTrpghh0lMsTdxAcr25E
qLcd/D+1JdZEujqZ+Qmp5wCoIV8bUZiX0AiePKpGrlNGOw44+SBNqEhVGcQV4bKc
fFqmvnix/j1ags30CazokraHCKF3TRzXdS3SweSUjnonqiL3yeJdl7oPVb+k5WKq
2UBT3t7SdQmIqtEzRrN03zNZfRK/u+kAgAQg1XNyCAvFN1npn6EruTiksIqkx4Gh
Byud6kMTrH7fvitLgyevCWnfxosgcjdUjsduRisnKz84Qm4KSiYiWi8AQQqSAno/
DKWtBi5JSgq4mRgVoKYMKkt8OrZH0zm0wpHzOvGnFVeRl6I/nCmAS3ZnkCLDXScR
Z+/D5SxnENmFRhCFk3A71dRUoYeHg6Ev/GVYvFE7byCYYV8wZjSpoQ8VyMnQXikz
CqHGpWvmbHOq8oeW+KQ8hP2vLLFKoPjMZ47nnzz6mo7P3fJxDkCwX30drvK0FQ7H
55U9RA6nV+J74IKHa64/Kiykskz+ECBmWwbOpwLfYRG3UqF6l8s38Lw7Dr4tzCea
rxjv5MJW1pv9Zy6lmwNAOYKFzBtKZf7/xpNKfzkRuSlOot/4/z32H3fAAMMr3EWm
ZSnrygeIapmOKcSkm1eLxQqnCHJR3KKRJ5VF2mJ2lmD46BHOwOAmXbrRFJZqjijE
OdWKUvysr3dDODmvBlPcEF/TGjlXoJqFmajkw6654A34BHx2+S8lTBNRHhgAv4ik
YZ/qvFqg+lvuXeTmUguThtl4fOsQKVcG2+ud0S9KtqjdVGdWuv/E1PZ6Fu/uioMj
fi9oID8wDoa6xxora8cCwm7vumF0hwFwkFIeSIes9N/5x5J65ep0NVXx8LkZ15Bv
X6TJwIgiVuTA/E1ciVGBFwtp2YT33p+ugLVYthcpooK80U9/kPqHjtdqIp7CpJcC
odPTpjjWFcLe53ofMS3dlYMNBM916ph/hcuNofZHLDKdA9nJ4g4AJyjktOqbYCqQ
VQAJwbj6QNHCuNqYPY12wZ1i7r3Qs0Um9xu1M7ocd91oErD3K5zyLtS+ZjTPmjZM
g8A9OvVFGbuOk3dLPnP3bOyQe/MjEYBqfNIk/Tjw1K3ImpcgLKOMLDBi+w2JVfyY
95LopFkVv93nxB7XC+J1WHJzg+B72rlRbkBlK6wFb36KJ66XNWn4Z5oXPOPJ0Xut
8+izM93kZu4olSEi+tKQG1w1HiD+6FMtBh3y0iZKKC4xWJ8MBimbYmcW19fxVAtu
kNi7IdET6pq8/7X2J24E82ZUgselSPzBOiO+7gD6gXGigwguoLXPS9ivvL05gMZk
E2v/oAW9W6kbO8gm2A2bkqpno63KiiOyUAJ8VCKjApnC/MUQ2NnT03qt8W51pPSF
1XAlnIKG1Tfz2V4JggbMrAPU5bpTUyOcFFbU8eV2jRPRM9CtWqsF5wKeI8Jfspzo
TW+rG/GMbSOaDtXK7wUKA+96NXCn6418LbZ3VWBq+RZxESoyfjgnRZb4yfMSC6SE
TjCUmj9HTVVXJ9x+i1XlODNJSvJ4bHh2SpO6TfeWEs2PiqmefMNQkL4WMwDCYQE/
aNTQPPqtqUx+2AHXi32V6AfSKLLSKquYpUb0SSNhs5vX1cXemNFstaIt9qLoYQL3
LeFL6GLLz4QB6lEKoUCXDO39C9K0m2vFBmc0AkLwC6wUBzUJ9G9nXxDU130E3Ssp
28QwsgFN+1RPEn2S6EOyrmplXxlkEUdXH5jJpYlSeJAqnru8u5eUmjFD6V13jxk2
/PilvH3GucF1bCiVJYaFlzih3gkuvv4aHd4yFPcUZlQrf1sx11191SjWkLb5tbID
b/dGlQUdK/kWy1JXDQZwzRpb/s7RjK+ZEoRrvh0RAf13Wa14RJ2nvTl0qZbDAdtf
HeS3kBlQw5uMZ5y3/STmSTnpKq2Wd9H6jTFsUbmoYDX7OCWkn/zf1ugHjfhoT0xI
vee6dbFWPKZIzPvlI9AOqP33vY/FNw4eNrQZRWbcotmkjEAzXodRSkyJawUDb8ec
1jI3XqM7VW6HNueABA9iuuA3dtpxDw5G/bS8q/Xp8RA9VME998nLuzQdgYqsRDn1
0l/Y5Bi+pqau7f+YZP+G4NFTFlpbXtCHW9Fk/V+FtPhpV6lEZKt9RiHbDi/9V7NR
BjI6taqiL5nM3fOL8XXufXj4HzXNygDDyctYW8RoldJ0XHfIV7PXyjOvOp/EEJvN
xL6V1qlfKWLaM7RkSwdFmcEdqr6oAnyja3LX9mwSfHPW4xNG34FdXFkXLvHj9bY7
pf+b73Kqq1NUE+Zeqypu22Ofc5rCdIGdZBKOP3ExcWzXo+EuFASCMkki0UCkg6o/
W4pjSpv91Vm7NKDoX9/jFK9I45AQFGucPYoq/j6uta3HNUOu6uxha3SlxY2bs8cj
zxVU3EyR/5J1ND4JklJWEWuHhHru9tvNOdxz+d0VneOF9A1m6rBbdcg6W54m41p4
CSijAnh1DqmpIDRs5fNhLkz5P8VtZ3XU4LssiOs7ZzD8+NiBluwEd9SYvgiGoo6y
0UARHoc2+hIeVfF+TGYHTN4dwCfY/MpbIgQmTmfSjsScDV94KYP/l48XXGczReid
61vEYwS7MRUaO/TfgUaJBzArnTD4mw2PgouDShP1anminmaU+iK9NNfKo4iuNFis
CCAurzzsqM2I/DtOB+crtAnOBrSvbrv66adBeVZECVDLKPIxbekkXXLkAUD42nPH
7Sl3DNryxonEHJMIroXYxUZnnzef5nADyHzTF9MdfqOa7NO4OM8EPmRx5dSv+J2/
gO0FxItCc0a046Z+rwLu5jgJob/a7GliDFqUuWYL9jSOjZr3gGuRA0ch1yqVn/+Y
0NrE7brdkr3jnMJ1/WfUroaBnxlfQqpsMeFc60xaUU+cwYK5ccwCK+QZEzb0ijQ+
WeMIcpCv6/Izsd8FdsD6m9/0adLRlX+3L6avMZPJCyIsWlS9E0gDCqDPpXVjAHdA
B+DUib57g54Y/Ttc4rGU6xrYma9bV0/Av32LF8j4aG3Q+Qd0lSIhmzFv4KWK3Cqk
Su1rkzVaMyfQOVhg2VGw/dPdEwkPnOl9TejFy/QfMxBoEIJh3JpuzTrU7Ukb7QV9
Jkbgy/X/N6ZCBhnVjg7ghiUhIscpyrA9FKb+J8QU5iCsR8Udj8JOs5HcqY0JnIKG
p+gWRukJgf14FvvCy1xo8OdD0WMtBM69vGdR9e+wmTIdJEnZ+L/SA0sotXFoQxxB
FrbwjkdYIOZwKkE8yFVocA6wxQJ/bKTHEvkJaJs4TD5Noh06jmw3kDGMvRJxWMI7
nRSF1k0xkQduoN5Vvk8uDSy+0P0Pb4KQkZ5u6y5E3Pm6l28lksonQQQa440amjfc
+JTe51thMzU6Ddy5FYkYO08pqlHa1KLo3b3ehqzex9kquR7jsvlpS77onhpkC2EO
cLFihmZZS+osrKw1d1cgVV4+TyXtrES8JMD3S17T43uERaK2fomtiwxAm2EbtIF6
+C604IySpz7bdSGhkvxG9XduTh5fEVyBG6KbTupwEbv7hPKnaxsk4IXcy3hnvvmz
3Q2uT1bFh6Y4tp2teg9CtRz7z237AJEAa6STbGVxVZYZZQtcMR1/SxZnNb8XqBdW
5CvFJPIbPe+cHquFUe4UFzpc27BfvidEICj7epg1cfiOFgCzjmuudHRbDcuX6Pwz
fUdhRzYRQ/OCDDDJ5ZUAqL8jyDfpzHG9pNx0PP6vFWlwE679xfH7q2WAGXro7ntP
afZDIfx5zrZvpEetPMfqqgbJcasPwW1xdiCsXZNCMTeGKtJY9825/S4rxa2ml47f
4wyCfu7SD37wxVZMFDBLtsICqcRnQCRPf9kbqI8wjHXZ+SChPrRPMf4g8utIxMGr
bltlQ254Oy+X7HBPu3sr/VtLLnnv6aZKqM/YC1mzcQhzIzrNt/YO4+qQTWib720F
qwMAKUV5r3OTRyAGKTEpTOK98CSSN2Gv2IR4lwNqk+g3jDOOwSlNLMWgZy+n5hpq
mEGDLYulV3iZYy9hmubcB3zK1kLq5vOLb+2oTytF+ZO0DsbXMpsNu/APxSAnS0+3
nI4pNPzE+BG4M3oacYu2mvgikpqS3v+rP89bldTvEVuk1x4NdBRET1cHAKJFY1Kw
l6y9pGDl4eTqQSLHxkM9873sfK+MPVHcPoojx88kIfjJ71TDcE4uxWmhCzlPFYSk
q2tiUn5uNualIdtRy564kTuAY+PtY34bPQrpJY4ZBuPX2WddonA/9HOaNKqchrh0
9h9DcaIOBjzK174o9MyY8FaLsafG2Hkvz0WGTcX/6BCe1HvWMT46vYdoJX4qHQoc
eEiqmceMjI0FJpniC+scX7C1+qakSf6NNwBH+O+NyMC0ibchrljFC1yrBP9tG0Vk
eCiupANzf92c0DGLRV4ayhwEt0G/Z1QpetAkNz7SiV7YIA8btJuaiNDrPgUHJKFs
pL93Z9Ap2SJjrgoTcZ5/ENkSzYB2YkJq6GxgFsUGn0MJ8YSSkoUXmWrE5GMwoXmz
4fg8TWu6/MHtiHPWue3suInmEHzcpv3BrPNYwEYuwMF6UsyOCbMybfz34UbmW3NY
0zqtadVhEqoff/L8uMI9GYhv+6jzIRz93NTfc8L9FFdI1H7NmfMrN5CZdWBsmB/D
jQWUu6FC50sgyarTYpCYQh0fJuhDMEvKiM1IYsMBD+psBknRFaA1bzdq1//VzXWx
4gn30o+T9itzXM0xEfBO5ScY1+zZ/dfgV1suIWa6SEtAaA+ly8OIhQ5paZj+EbKy
MRaqKjzExw6IZDoOTwXrs/J4y7NhkaAanOBjPVlRZQjBoVSjhGclpn/wHdFnF28b
pdK/JBBEhrwXOZd8dfr1hRD5dgpbF5SItkImcnOkxArc5439IBdfPy4dbIe86M96
z3eZU/oQbOT2dcBqzQHicSYRJFGzMD6k2X2nKdsrsDTxBDJPopeXZdGp8S5OTVM/
6GnlVGFiHadp8QVoyDNx7N3GzupdVhHWGKc0M6jpcD2FK8DRP4mjEXMU/ji1ahZa
Dyl8rLPKHOIvO4/AXHBcjpo12G6O+zWQ2A0o6HGKgVc4LFR7qZzsw6zSDyUkKXM9
KsVHB4YBXnO5+mnyxD8XSSK3Yf6Isp7OQuzb6DurI8E+uXAd9wlxh9QDqPPJ3/mG
uK2OLDPNDNZvKX4q7cuGEeHdTTAlXRNJIFrjjB4AdOmZQhGQ6Z0VtucFo9zCkWZ3
g/FRSiZGKBF/bXTEVL80J5pZMZr2p+XgMeVcarT1UQOnFUj9rXy/NYGEdCAV6R4N
aGTIPJjMNm9GHDbzju+zXFABMw4h37fPI9erRv464ZR3FjIfeRV1YxCwh7LTSggm
/8vheNGc6gxclp9HwabASDC6nTHEVdFtruVKTDOxf5HifhZuLKZWQj8Emshcu+Z/
mmCBWU4MjzCPWw4w5ebVivBiBf0DVPcKw1hQ5GF+cBTj9dObGbui43igcXDbB7tf
GkX84fXsqzFQgeltrJ0ENeFODpOLH7JuNl9crrvlouA9A1yYZEjkqqHefVJ8B3N2
fl/RIyAq3d4uN40sHAOiBPKPNPyCAdFk2Cs2SSY7h3j7JluQDXVAwyF+EbJHDVLU
yljLLAhMOR33MCYvgX57jeiQLdxeGH1H/W7n68wF9GjvJOQcHmapdftLxGSYIZKK
BhsWOjj1CZpzivkGiKVPMU8eSHs5IDC2IOlJEkwXrPNu8w52DhSAgYwxUdpPLcHy
AcrZwTA7y+1HHp3VmgSdISm4i3XBC2MagCQ3ntcfh21QYNVZr+sTlPfqbXLVvtH8
8Q7e/VTW15DPqHKzDmoDH9RT8nfIEzupChbZNGHWw1+N4gzcHzCBuokQWyJtG5kd
AcdsolD33rbqc+ebytG2ev03Lv9kjD1OZsdKvfBlePsP7eTCNr7r2GXVm5bAyoN3
9nA1OyJ8XoxCJM4ad8ViP4Keef1ApmJjZOiXbAlXWNNNqM9Mdyd0Z1VlwZ9Lsj9P
+nLVwde7L4KoJJzjUY7HMxFPlMWx2ZLZZUfaQNRJXy/pxXJSkTF2FZbpNEdzQGlL
5mHeNFDbXwpJ6k3flkRH4v9FRVhdeSZkkaiouuorDF9F6tfWOEVt2c8C4SytSEPY
r2zFHlhPJBtYgBPTPxU4NApfpIaaEoUrqJPZ6+lAjMXHb5B1yXC+PGp+2AVyIwzp
kYKASF0CGbmx3U+8Tj7S243p6zMGFYa0j1B0ao7G4tBmD38jhG8qjEWk0SqBOvbs
LiJJEiCUIVxiK5y8HE6uIQBHxZ2XXCH6b6AaObJRr+DeIztLA8VDGxl9w0G8ATyd
6drf1RlaDwc8VyKb9RGBXUoClT9efr2zsqGxejfFN57c559KO9Z1USRRlmM0Gt/+
YZFeVo2owXL01/1JtQqyFCxHmToMDORTlst2oWELmA+SpWkvhfzoRK2VlwLsurX1
Si2J1KvvUbXPTrYFXsdt0nWKCqn8Cet1wccvFWAD516LXCIZUeWsWOD1k4KzsXGS
3dqrtmaguh9UbcmQqFQ+cUDX4Avmcb7XGyhAHb/riIyX+EuFYPJJ9pPdTJSg4qA1
+0byJTBIVlPN9E9EPhwVeBNvewtNa9mvXgcxzASCdD0emBjosJJ/3H/GF2KsIYie
9FvTARLNRoEMTIqB1ptWWjrEqalR1a/g6NTG3qpHjtf3e5gcBzyMYO9fbloS3UVm
mT5ZpxU0GIpcHVUUGm7jAqOgUs1m06FMjZZIzYC7kiZtem4jl4XUGl8Z641FdbxI
SmguQwUf38G73ypjkssNWuyYT/LrxMN6IQ5lCccEHG5mJZ+oBXMblnZ2t0A1sQC/
qxOJE00toQTdMYe9Dg3YtNPJYoocNOHUiU1IZq2SHfPUM+kMaxkwz4kqcvJ7zCrc
rU9SPM9Qo0Y+8htKMdCGdrjHdth63TAjygXBIlTLu1hTVpfHUYxyVhQvXLlKuAKV
EVKWOi77xP1H2jLuZKK/kgoRhaDKXZPEa8LQ8/UZ1um2YKejSuHWTAHR43TKjtxr
m2AOkg0h3t9zi8hHTohkKNcwdw2zZBarL1tN//yJ7ZHWqekDqrV8WQeRyOZjsquj
k7w8Ux6/cNOs4YzOGoO5uN4RVEqxrwMIU06/x1CrQ1E7LG9k8fU52zyqG+A8TQgR
WrL5SMYmlC5qQowbzi4f6J2xxpKfpRcApyEsHhpQB0UjSTondzEpmgAdOFIbh9oG
pQUJxbJsNqdYYl9/9uB5MLTzz/i/cRljVUVWHlWiN5qdGi/uecXvmE3O/23q684p
9Txe2ZfRAAdg+7CdWfDTPoLhEPJUZO91ulfCafC2JSyOO4XM6qshxCKdIOhrwGor
dfbrosky/4T01xsao1wy3IOabjfx5/ZDkdmGwVxmIWCiDKyHsef806GtBDMfZ3Kn
zIYcxudDsro8/rPDrMrqkt/c4VHKNAro07A6VAwDwMY2e2T3P4Xitpl8dUptlCt8
SMFn6gRBOewuOLTlzmh77OJT4obzKUekJpuwBLpT2O8Jd3Z7bDWGB8Z/l8zW873H
fVef45sH11GuiLKhHeLlb1xE8y+9NIIxv7Nf62hXdgoVQQiokKwunxQ/QxqSooYC
Z1WtWvnTra4kDP2DwEC7+Whf9V1UafLtYwOi/9eHXuGADaoEKIQTF7UzU6CwXMvR
oj+8WlMAY9A6kO9t0ZyxnbMa03h68yXeWrVR6xK/TradSqoqPsXJDKYlLZvv9Zh8
srWcwtu+5gWTVbcG+RYOMUIsTZLj5AZOoVdup956r/wWxODa4UfxHaN8B/Gg9UBx
rjZ9P6v0jHKRnIuZVeM8H3deKqR/Lk5tf41YF6bRiTFhC2zF5mylQYR7VHsMy+FG
KXtlhQM+sYBp3KettXcsjANZ3l1usGZ1bJ0rVGA4IxOQIB/xdzTxYlK4l1xDtfAz
oOi+7fsigxg08uAvree8tMroqjjiHNbfn1KP3K7gFW6rXiBIi9VrsmTKgFPNvuI7
a79ufVLZEbp+riqAxKlpoPF1hy3ElWzsgf6QC9iifivv4MM5jSKR69ODgmAVVY9l
BD/dIfmHfV5Qho6d/oBrX/Khs9e0L6+O6po52shFpJDMwJ73kXlQylLFOIKGd21P
/GnIDnHuUGHH9kCr1PMoRcs2fo2XofBtrtjO31fnsPMclPm6PqDnO0fGycq3duOQ
9cY+LXNkUupUtfYQjZKOAHQo77/SP3QsM7Cjads1aEYJ8I1gWAAjHNOkvqXXhpIf
x5FyPlY8M3GbVeXKBSBrpeMsa17TTcBNW5Xsp7/a/slKN5VVh+hvFuv7xJ6eG/hv
LXXIzW10jA3E1tezir+zff2tL530QZgU1s2kDXbEA4d3CHpUp3g6GuypotpdEGj8
jc5zqQ6B8jQzLLC302Tb1vq4XAGRqJJWHmpju9bOLDs24JyOAL86zbg/U/4+Akhq
MlqxqKTr8sBuaogupc/gfH84bu+yczrEbj4QC0kNbE/RD9QegTowPsP7zYU5R3Ot
H7kFrlk7b42T45M+QBRUdsO/EEOwFhzR19tocd2Gpym4OWBGHOND+kXoeFyayBxm
heTaq9kicDycqPvgJYwD1XVmtBc9Yz/gtUQ0F0C2nNgsfEGP90voi4C47vNfr2qu
mEb27NwjMnuEHUnwT02gFye8oKTQUjztgjVA7uowJSwCJvUNMhx+uSygssReoTn9
44eYNJWGvlsVhDWF8k59DOVATBfZWurITpSwd5CXi3g3sKKi33RuElMicqdIHr6n
YNBKLX3mrLjWyJKnN55Tmc7PTZXYHB/u7s5s553qHdJF/Yil8gajEOWrxp79C46U
1vdAw02K8IP2Wfgs687LSkrod5BKb1DqfMa4y0ZkMr8CG7byFtlt7ssC8L7E701Y
v+MoFbtg3M9AssVOsPEjU+HJyQci5/gn2S4GEP5nM5a50QX51C8T73WbRSfCh9N9
RAutUfpHKw08DYluniiMHG23/indKnX3LYfH+3UjjkXKFbIaGnri2PQSwXzfwnyH
6HCUfxv6V8j6UrOiYshcKnrM2h0OZZpX094EH+I2fZKJ9X9iIQ1XdfC16dsXQHjN
b97+JnEjxrCYEdb77LpEbVmVbqmvw0HFz67zfTaC91fJybjSZbHmmFKO7w4r14mO
rAyyyPrVUQU6XW0XSCnL0eSz+StroulX9g2L/qge+rXyUMngtrOQOwcfjp8/8FzX
C5lc/OcsLVBz2lUEo9jUrAs7GqXnmHkWfCohS3Ki/dURBn3H78bF13SfV8tS8vvi
D02T5xEqyjGT5ttM1VE8uGLSug4TinIhumWHpR3Rq0gnOiJOL5gj6PchlRF9orHF
M1tItn8z1qHcG8odI+MRI8BJk7G7SvIXOhU/Ik5MXZm20RV4NWnb4FpSAJL5PSRu
TLzbkYF0XJISigXtz04g6RmDulH/LiJTx71Z7wNIFkq1HR+TQ7LrgtAXkdSkID1v
c17FIPPEAfPeOTQo8afVNFyKZOIDRHTb9H5+e4Jo19WHde/49o83Lky+5BW6+Zy4
yxc/wLN4n/yRbJiIFS0wFNSZYzGjspJUazMaqbAqqW2E7Bh6n/hYbHqefq8+JQl2
oyFI4+Kwe2YpKHLqeSkuOiWkkTAx1E7+aqUGnlRv+068bOTqLZ0SjgyppPJcWwsc
vfl2iVxPg5Ekosc/VUBuSNK7gHQhyWTyI8X3JNXT6OD0a7q3yRcnv8RYzBC3++Lp
COIQmSJ1uouBABFf2c5wkNp2qM/Ft7wT1Wb+/qwibsKhqPIHVq8uAnDYaQpORqs1
3jMnaq7pZqKL/HI5WW4g1Xdzv8BhDfu/U3Tj6MyU5BIeC0BxRmPY/2tskG4dWo1c
hSsrJE6hK6VL5e/wfAR7Xs0noCdgz5Yc3ET7PwCrHa8fLyGDwqvXFFmNy4lIn2Xg
0H+nMhyf2+8QCw26tqbUz/c/YDQDzx5bZeMh3AbD3zaXfI44vhcIMTvPDvNscUQU
ref99DnhvPWkLHXSkBF0jJQWtt9eaDmcn30BSbY91qPZXCp3jcQ2ZjcWaWFUCqbD
1P+REHZpJPUNancO9qRheXg/BMZVnqMy8x04+OubDe9g4k3Ae6MyOJqlEwijCdTz
ACBwpzE+y6ghNsdj3kDJ/KPs65AUnL0EVg64D3sdtXxYQyQXee+dOfT8o9hFyr7y
XmuJE2lF+xD0ELsHAm7eWB5Ukc9Zi65RW7FkVu1SVXVL0tA2OcRS9kLLoOu+6Hcf
ii5p7AlXYASGcrCMUFGrajeaYcYvDyvlYkgaxcMrWPSH7FuBIfkitXf04tv99RkH
q5YdDweLRwBxxUQqWAAAPO8oyswl1g2a+yPVkqkpI0f2Jnz6lF+XwSSQO2pTqsNT
SWDU5QH/OvgpTioqD6KvBQa3lxBfPZbBGj5KO92J9Bsp0JKO6vaD3Gv0Ph1DiKs0
LvvJt/ZdF9QWD9EtqY1VgSj1XzEwk73VZjaJlpx/c8scVsDODqlbh67UMTNLm7/q
GyG8EleKbJz8YzrZzrWtfqexNjYkez1hiUxSEUAmencEgYtwxslI5qM/M14Bj6ZX
Q8bSNVo0jxz4WgyzJ1VsZGZ9y1pAPsNY4CM3CvNGWGuSDUWBh29w5rey/XaiLpUA
lC+JsptS0Pv2hIwt0HVud5Su2e2xi0ScFyo1qp1iM4duJJgf8o+RPjz5QiYZFM1p
vNF9mBs52969aFlX4eGAUTmpwJytvToQvu7trcFfashe8vmVvE15nBPvA99x7sP9
E9m7CcB5xaf9/2XWfGYx/Zb/AdZAvoRy/PZeQA7gE8+cJAQlb9+cADac/3Qfay6F
iM0k+oapK3qr0efFhsshFWzxVWqLD83PBluZdfo8NQOHxF5wIOuknbtq63bbI7oA
54WOIIlNFwruRKwaXkcRUB5JftYFw9SSP2oxUbtRbXtwt//qpnTZRcQtwD0dBq1J
cPJKdvv6oSelo/TQhDL5HFpNJ7YdWSNp0Ozra5PmsbVJy970X4gdA6+3Mkm1ONMG
lwhULdrMh0fIRpXkWMIDVddiErx6cI96wdMdeQzDIKS3HKmXdyukzE1hhKOrL8Ah
bDYu+8GXZoYkt399i7RDiym75VymoE6zBDa7v4hPg5bo84Lyzp4rJcCO5yfT7QsR
CgPm4lAzJzdmJn6h6b44oSgWuk62orD6Qb+iKIKL1eoFB4VFunRk957tbV8GSTxS
L6BJruGNxGe6cSjcpXYoZz+8ozat+EQYN+Iyd9GEla4xYVAJeGRTlMEjtNO/EnlV
RizCPU1B2G6Q7/snQc9JUBjfjWIfU0iL3tuXYogAQArnEFpTkAT+oZD7nMFGl2EA
bPCfURIi0TXlApHpwXg5KcwvHxSWbooL1Z23cUPoWmSlAVcT2Isv25/ChnlSC/3K
NsBhvWm6SD3Q2vBiRC3hQ9lv3pawFoOSm7k+RwAopcgK5ML3QipDcJdhf8uzcTYr
3NqJKbMCiPFp0dg3NH8SI3/HZJW10lVsgs+PZBL2LjS8/IMZLM44KM86I8QufqrI
5oBTLPiZ3wvM4iniL9cd7+GQPwQ9d8fBGaP+coSkeEgV6wLflw0LEgZMaGx8Ee8H
N50xqCcPlQVrVT8LbiPaWYFJMVgb7BlRzl8b+3qSCKumdvKynjw1lT0RBIQq2fEY
EK5IIdoBURLMG7qsKKUVNLvgiRfLAsecwDSJYVpHWDBoG8vpFAq4kZUwAL0eG+uH
i5pI++THfH5qan8qbiW5jaXlk1jsEoRIg8uEDd6/FmZ7rcEwpSCfgl1kyrAAHVF2
lSxU5s1Go4ehnxhHpGS+xJJXWEyuT8d1HlLwz95ecExyy4CSYHEDYfW7MdEPxREY
hujuPkpZnOkzIie/7EHDdjL+co4DvGbcE/P/Uq1WdjiU2hQz8FpuA77e7Yr41NJY
sMhMl6DWEU+92w4fwvoSeZdriZcqmDnTXJWqXRmzTu5fFvw4w61Gtzk2WvDlgwux
YXNd9xPFHooqPDXNsiiopJNBUKba0eC8kewP8r9yUTWVEI8gcrLNvd3BKVFTH1Jk
jCci4T2vI08wb6J1FH5VBdDbEWNFSv5+OqpMrsY2vSmNcFi1nL0Xi8R4MlSpi1T0
aiHk7bp8B5Bvp1Ob+t4rdOlBEJfIbgG4fGErtzgNz51b9QmhRE7FzXi1pEXLL97Q
irgI8QxktWPtZxf6vuqq8nirKEg04vZvUDPNb7+EnFpiwIxVg+zDYDVasEzLk1pH
gdy/EDCvKeN7Wo4274Jeyu1ia9x7Jdej58cG2pzNFXOnA4WTbiFcFHBCboCrfXLK
TpIXxpWfx9YTy/rJjskjxBTPegYxRXM/zsvcHXE7koaQ4A+DaCiBWDo1wd7zHEVl
NtKsMLcvSoRaggqLnuCUpTFo4Oi/gC5QPhNqys2xox4XcntL3+CzRJ78z0Csmo7Z
55kgi5lcIdM9UNB+KeNqJgFvO9HKaCRx8QyTT+gS6ZAQFgjdzHuAcDF4O/o5FSw6
cYWEydXGycV5f62tHWrI/Ex9D/jdblpeIqkI1It5U8yieChsRB5xCWs2z25GCW2J
nacX2iQTPiMBNYGsd5WgZjkbwRkqhLvzUfPhN1t8+4G/fWuBbpkovmF7CoJJs0ua
KkUJyS++LAcEorJ/tUFXJvy1kK9H4kOagOBWe5pQKSUHYzs1dSK7GtSEvpZ4SsgX
0WlklXgh88312oGTgDIjirjamxLMIfVbOLuvJxdploI8o8NfhQ20UUrmnTeWemZ4
7F+MrKMwUvMjC5Y06hyugJxv9oqEsCKXgcTQx/yWXBNwqYw7TXustY3Mq5DBLQQD
L8zsqXcO5IELvvkd71QspJRVIMXRXdbuK9qWRMAtfzWtk6QuCfCEP0cyEDxl+p6r
nDeXbgkGVvMwKsU/qcEllM/SGX/83B1a06C7BtXUg0nvkCB0HgHMEMiLVGLKvTHF
V+ZSjezuGXS0ANdQFEf10XapYsP3TLnri946D0XNEscQ9mg1kgkpfvG0kCOreSN4
fy3VSK1IC/OaDakfbEvAazWVqc/I4hPAbS77+tlx8g5mrAZVGL2eTrG1F5aqw6AV
ikUmJlTz7ECtjJjXi+5FxfZk8qy1aoz1k5xydLxYsGe+KjNK2laJiv+hPP0YrNJU
sY31lGKf49GLjnqh5DeSfXgdpkeQjfm81onYPcvKjHyHK+v8T9kQC5GaW8n90CSW
q+gPuMvnU/dDlkty6ZpoQ5YWAkj+atRqKlIeYX8QnAB3/+P69EddU4mHjW3m11H/
aaYu8sOnU+oOGtv4JmwIEF4DxSEi3lT/0/H7ZZ3bzvIGzGzwkrVhZfYK6HWc126F
YeMKcjuTLT3NHe307kVK3dYvp7K9HaOgWJvhqo5ISruBI7e8XXuA38ptAUZ/d0C2
Pxxw0h7kgBh4g2Q2PF0aaErB1Z1QcGcm+iCEDmqyDfWy/SX6VNAmfdOUOix2dmn1
AYRBXlO0rXxwNjSk3kNF0lQOD96F22xzlCOGbuL9DaI/6nF1oMRY1OyncHqtIbiL
4zJ8QVWQjxtrODNKieviNVvLtzW+F4Oubm/8JKhniMYLzmI3IY9NG/h6rH3JRFFD
fZy8wV+pwAEmeDGdhDyMouGNubv0Fw2BROiEeXrpWg2eYDlfV5BT0BIEAnu2wNSu
VuClk7d+Ocu7pdiBsLo/KlZzkZj2AOjS6F2sDNTzoJolkZoCp+zlM5iitIPPGOMa
ytS8bUc+bYX+AbeBnrumNjvtQTYKoqKrP09E7v1yqAy91ru0H12df5AZrh7+YL1E
nN+GNEOVYrOYk1nsFQPf+i+MzcQ7k/N7DtmrtathYBkJrzhTPilx4XGdoibyvnAu
id58i884QaOF1Aptp53Iosi+9kObB9o1TY9mfYHHzcgvLfCztqbFuWCysn8VGosy
/fI2hqus+Jr6Dqfu9MsewnVfthvwAuE9gvTKraIqz3Rh1QAe7YJITLe1+5KXtxs5
XV2gPgWogDUbn6fhAmhdX6ABfgU+CJsNOrvpR9snlHYsHgKb0H7KVumgRtOEoYkO
LITzBGrEpova9X5w3HS3/8ZuPYzaYzVtA4STQtonK0tOqtz+4qVz39FEon6KBKLj
AdMaN5Ki6ssKK+lPRJTD8VKLS1L9xmgZznxOnmXZXNHjXRWUIdfCWZbl5hOpsOoL
Z3LgmkfIDJ5SYW+JvrQLJZpUpaltVG4Cmu6RUkmtN9bCRFzPy/hdLWbHofI9+1ob
SYxFXfPInPku/+bMmMK5qLPuBn6cqRubqDVNm26ULvs00HombawrPllVa5s2ZWgS
13TA0JzspEamsFYKUZkM2w8Mg0FI/Nn5j4T5A+0rk4SmWfWPfYCQX9plHMhrwRNz
3L6mQ2iKl98eQUHGZgTUTl9kY1oSeZQZu6Y5LvGbIXkdvjk5K8fkaVi9OC/d/Fig
AgzzNUg5dIwUYbtAs/CDm264w0PwYrEp6czdvbeVRJ6YPUXqtKBm7UHlbMoFieLZ
6QgjOcKWuxCpv/VSqt8AMYwkkI3TYQKuurD6E9UR3paUxjpRcrctPG1YNwn61PRx
Vb1QkmzxTan3pHSwIWC6eQeSx6lTIX5h01/icx3bSdyMKc48U9cJFGlI7W/7LaTu
2PPWFi6Yxjl0a3b7ePn16mg5j8Qk1gxq+HVZEeqYpJrTduzu/u0uSScnwk55FXyf
AQOipsbJ7vltZIEYBflua+T67YHFxy4ksEAKlOy26JWSRg9ljh92M4IGqBywFdo6
6mN8g3bRPzUWNYfb97UnGNgWWRX/IJiSgth53uEe+cbqvOWRZLyqHcjAEA0L0X0B
EWHGRHJUl6UXi2UqMmZ0X3mScJ5aMiW2pjh77zDJ6b86uqf2FspHC2QPEtvLLQzY
3fHsO2kGHGZ6L/Q78vrkfCO43w6oSsDWgZsAsTzdfRXvGrn1rGfbA87OhoCRyJJO
qJtzRDi7MkhG0tLojTbn51NFk8KN79hxB9oE5y11GQNSfMawZiqPPXuty7DYw22f
6VWHeiR50G78u+PenxqjYpqZM+jRKUdZc7XmZekxtf7970A8NwC+jrJKc8NnpXT+
QEvkAURf3QhxYUBAtJNhWxybBEcobLV7lm5Q7TOcKnXANW23MIJ1nuTzZwx6F5rs
/sBF3m5tdofT5JXwlDQ8JPmekM90U9BWADXLp7SGEUQoI6XVs9WSyb6DNrwgunu0
9HRt07SANSHkfueZxHk5OFtCht8xyzi5pxMYtxbHBavw7JclRokY4Eo2TTOk5Maq
xmMi5sazrnX/c867KNFRXKoHliAzBRAPeXLY/4myk4eZ3rNCtQ56ysxnvd4PG4uP
FUsmnAsjjAI7F6ysQDjGuWgR++gK3gmCDt0Pxl91rd/J/Ml0z683YtdOTGxREf34
hMgg1b5ss1i+5Pf1oHdnfYTCavNumgsGcpsv9gf6JtYHcbs0Lp2LRvp44UpgwhRe
TLsR5ttVE64i1XCqdd8a9ZgTlFAKRGm7wgf2dzYNIJVAEROZ8zzLozMhpfo7d2eK
c6keRkBbGrRJFLjiqoCP7XL5bN5MXlwC51awYYvLMU/lSCmDE+YB+k8LH1bM8T5n
F+Vy/n/vf+UxFCea7VKOCbCLpO6YfKVUEshSuprOBxQl3kWe7tHRt+NbHfi9LktZ
ZS01/WCsLg3TkTrIn2dvNWbxySVMykaKK4lsJPdUzK7bn+J8h2JmMNIW4xAvnVxe
bp/aVIEcr9XExXgfZBJVFOabIM7R68AcRnzvKSH2leiDplbvrxW5btmvtIRd3AbJ
zsPTL2Ygol49o9zH198unSwHxdgo2bcUPFAgBzwQbz2qnTVLsIFIpdZNAvK//tF9
qvmnheRIBGF6UMK8VhPBnr6/ktHPL5zZhSVsVP8bDALEDYrk+DlCWb/L96Ykv2rz
sfvaUoaIpUF9o77KNti4PxUN5/ODSlCJoqimXVmOmSyIxxPNr7mD8Azor/5Gj2x5
74QZnEybP5nCsT7P7p6vBAJYbCVKPZQEB4Lxob1GPuM00mq92SGkh/4cWknup0LO
YeoiZm9W+FllQ/EnDMrn5FPzGCbeDHBqZInE54rBJGTFlD5EHnIaqwrNMeTXLDJr
Axtpy4WXbwu5J/xFRcMxIjcg0AqbRWvSDuIDjiLA9+lxLknjxGoiHjDswAp/r9Cc
144y0LMXQCK14Eu/NdolXlMXBljy9Ea4vM5eCJThxSfEW6RfZ7JQ0E3XbXxBHqYV
INI5oVatHozWMvmLkpHTdwEe4JTmkNT3yWWruFrAYcIvFMh3Dy0BlBe3lPNC9Z1S
eyIAH2vOOCPdHgsJTmUFujWey7bVkRqjbPo7jbEBQ2/kaFFDUC8AiDCFiAsFbCp/
7Q2BQhNMMZoYlpE5PrBMxWa8rdlonMqlgTUCriTV80D6bA97Mw8rH1bgs90t14dc
QmToHjNNC2t0RsBnigG+TwkePlLud9caKC4lcf5zdFeGARa5+pBNaGHntXln4D6Y
odbzAn7NxKzoStU0p8I9lrNbbEjpLBH94oKIQb9JDIKgn6N8M7s7oZACpnBl/6K8
GXL1MEUQ3GAvDt0OMdWxEFfQTMj1kzzHmo5cA3K48wbA/R2k9XrqlczIh2swIyKF
hhMXHntSKak9c5QeHdxND/AecuX+WPgeqPEE/rlxmdSg0bRB0dUzwDPcQo6v0vrQ
YJII6s/6OUviH1/q4sIIgvvQZdMJY162y2TEQEIg7+pMWb0T3blNZs+tiF58vlXW
y7gf1ysDv53liEITlMsoCzxuEPGZvVewC+hMU5OkxBui9jfiPRQuNta6mcrfhnSq
tIprQWJdbA3GD6fAM+4wSJo6b+Ol6pzjYfX+/SWFqGRk29OLR9ts+n10CqbIj7DZ
b0m43g9b69tT4OSatmKMpFAFhhIvuj3VJ/JwTLf/sM2T22l7HSVGohAtUM12jEj7
P9tZK4SwOgTUYtSl6AaWsMxh2YC8KGSKepQJcrfufGEZJuWyqlAHmgzsG0GncMSY
rsvK6MPPDXN555epkEQW0M1xFaf9ME16yY309+cm89elRZaEyCgUyYds1AZvufZj
MPcDFgvTCOE+aXw9IfGaTEjb7U9CCnFvqczw5cKyCACZGxQBWBepDD3tPsOqasHJ
ehFlwrTtD1qOhDTtEcE+T+3KFZ1fApyqXBtiTE0d14LcnMSxtsgLFN1OPCMx9RD2
xd4BKQMt1SoP8bPf7JqmIzWnXFyONqTjhbDNFQzp1PiEgRAE55rn950U9LSBa/2R
uP6+bC9fWV24jHfdUf/ppogLuxiwWYOPiFQqWQUsRf7M1gZpHrq3AEyCXK9RowgC
vZ+Djpaa0zFuNZGJ7PRESJ+vnHwCIU8hQfZ9mLty0LDQneErE6te4QmDOriYSIEa
Hr0hy7aDlLiZ0v3LfHnyKiiH0A5avCR5lgdCT76jCJ+ayB7yUq2wDg/WS/K1E9P5
bb5uPkdXzetey30SbXAL4d8Wk98hc0YnqWQPvhNItJdvxsjCgKMPH/tTFoFurI1s
QrbrleYN8Vu9wkbZ59Pv9y05QD+CDYOXCTuTrmii+RIWfDA+xwpC9gfbxn23yM8l
BC1TLFYiSViZzb735YJ4XDNyxSA+lObhz9CWhG+We22UPcanvJE8vsYK+q8vWe92
QztBFOFEQp3r7zW7UFqXtvrvXqlQydWOZ2eu9wDxLrfoLzh+3ccQuul5T4R+bn/w
jJEmIvIweQIrEMwRDOm124vVifY/8qx8opjmHZR1aS5MQealDvQPObXYPBP0XDXL
8J8FV2fwHh7W/0U8ffzQF7JYi6WNGIn6+1IFwOYFGjlu+n1mghqQUrOQyaeMw3Ii
d5DB3jg0tzRCuSL5l/hHoQepXe9ZVlQk+3bVEsPJmkToXrkdTVwFpZIGGhFIuW2O
I7du1Ra13qUbJWCXN52Cb1epTin5DYTIWGhcUMjmizWKGX+6ekGGEKwvgXJtedzK
gpe8ZStG5dKyDfwCU8Abihv09qH5MbDqr6TtOWyhKP/K4QqhgWgzJ2CSLD0SwuNI
j6ohWCwEoBI4+6odwO6puEXKEt8Kdd2DVk8WyFOczABZlXOoPglE9N78NHPJ8PRa
mT2upTMiNQ/RxjEAxVkd+DycFyD7QnsYC2fU9Js0RPPaijVck+AYaHK7UbQ3P/lY
x7v9+9YJIViF0Don4/9+OTWZL/SHpMBDTitRFcfnpwwMxE6EeiduHxPlu9oXKIk8
HzcMxihAPq4w3d7FB+AbK+k8bHsVoAkTclCVjDDEMMT2yYPewIfYVhesACSGVYpV
mUyL5KB6FDxsam6xwTNbktzCPmiFWTnzDo36EpEH+qpcbidfq2pDP2KcC4tjWc6q
c8BNy6qsI+HXx4BHpbzFG6QzsTcSVUxwxVofrUJh2zQ32VDBydbKKGwiWfwQnhO9
FptG/a40gwt4Yf+cghBPvVmXlju7qhfUlXr8ipbtBO9RJV7ENuEABsKBdAMVAEs1
ykA/HfIVQxv5yF3OKcDcxZM0mJ5Ow/Su2cjsf2sZfUKa0Iv6PdMSM6PBK+hYMdMl
kdQ04ju0te0txV48m7IxjxX1AgGSKK4/sQAvY6nfV9fs7pVjRBFh/jcKZJXSTBkr
NpDyawIgacOJAU9pkKI3Eh2Js23PagYHaUmWxhJMPDL5ZRWF+zsooKruZPaKo8J8
XtG5o4AyqkTv7dmPCPO34r6XGOG1auOSCqsPWpQbl3uBdW1vbcIY1prycQAqoBSK
XbLd7dNqwbPa0V4IILRUDL4f2dZImDSzGaKyfUYKlb0oflucWzVQOO1/oMYNbyoC
Qg5Jwe98m0AwjsdpSxKuEMcxsmAHB/iSt7n99zE5WhgZq8wAK8j+0VizMp5DEVPL
ZPPau+7sjQ9qyhsPMhq/HnExwEynlubUIRVCTEgNOlW8NjxvZ/4hJAECmaJisXY1
sBlH3cg4AuLKv8cnQHv7xNTo597XUtm7qY0YQHhw22Vs4Iqvfu+NI+BQBotivImw
PEsgjmpsxHmcbdhiRO3R9kof2SA1Dlp1cJjsU2KQabWiVU+oICfJx7VAJ/emcUOY
Atir715sAgvvNnpZcoUwXBpNFM378gR1KXOl24k65gYfCvgg2qDaORUXPnPOifU1
6g2Xer6pDh9w55d/IXOS7ZR45LrNqio2cFdfvgqG2ZpcN5euzHvaYsv8CbEshL6e
U/wvNgL0W+0ZfGFZWlyqGhUGpAuFaLUCtuNgpKYQj2M2B7RA1RBDkMX555S18tIY
LmJNqImL8SCu1AmyzwpW8o42KZAbRKVItvEzHu625xatI1UEigp3uzw9Gf2nuYuA
wffT6YzKSYEWiFJ7Ng2ek5KCVkI7MqRN+xGJmivl0JrArCHqPVe/CAA+XCDqp7Kb
fX69M4S8IUyAchF91SBaOvKUJf6qxDVKkcKTa3QxL1qJIwDkfDNL1CAd9b29VE1r
r+BDbwLX/CKX9ncyjrRoKz+4Wx+VJ3ib1bnjkrCSFXJO9fuFXyUXSEoFrVA/jYkv
yqjekaTl43S9p2tKKDyTcKfLV/zy9dm2JDSnc5RLpfSTBFEyrgrzMa6kie0TdiH9
BRTjcR7wf3IjtQ9fpMFWAPlmM0LK3rb050l0ZPSGIOq3edLOTpIV5z6nvQbQKVvN
86QZMC1+/Q5hOqVTWFSaj7gZPM+MwNXCabEb8yXLx3UmX9KsLzdgHbH3rn+Gz33k
VcUwtUxYSjvqGsAcaRSDP94Sr28n41dZVjQ69SKHJaKqvslPCTb7gLA34aSroT54
95tGU/QqQsfwdljjBbYgMHcMpd3Du2ZhgoDrwIGsxNT9FbKJoFqdeK7+ffBWDpeQ
mtFZZG2JSzNqD1ULaY+0s5aZA734tarciugAE5k+q/h7HmlTLB16jMfHR5/orbF1
Cqjr6yrTxYMnn1cdkw+QDikSo3WEZ5ogdub31J/MNmWGxXzMAhG5x5KEfp0lNQYR
clGrNTjVDCY8/9Y6tkIwjivyVhmzq2kDfJ+tKhpsWYsWH3Zp8RTg1vHJDbEpR9hg
WY+f1EkqL2UyCySx/5Wq2w1gGynSe1jczyTfTiYLIVmIcr36eP6lJ8XeX9NDSt0H
fDL1vrsuuzoAub7YbhcIiqmCiTSz0jW8BsPr2LecC3iscFMd19NsLq9iV+LaSdWX
QxqkFqqIAlPC0BAjzm7qSlGNBvirypG4w1PewwVsPDTOrApJZsEo33clLlirRskY
ezAn7LCXpyvrnQLPYEnYGyYIxaWIVpHsVzPhPfh3cRHIJ6LvMwHZLcEzV641nN7V
n+vMnA+kr3CKNRAA+wYb7twMeTi8W+5Ya2BcqtMfTe1LXFUvEyX2/4uHOGziY1gU
XArYu0K3S5FQJzIvCr5icoHUcxgTzmnci/l3Tn0Xav8LgE1MROFj/yznXDTnaUrH
H07XTm+a6u+db/VglqqJuHhL+oy1sB8CvgAEIZYlAEaj+x54Pc+COFUEM7INj9N9
E2Be95Vd513avE6IfCYB4EakTsEzmDboUWx+cLIduqA48jxazaCKWGpDmKLFGgj6
CPt0Em3ILxJEC0v9MSe+KN1d0qFGlVt48Y4YLGI+WRdEJIyqFKXHLwOSy7N2SsQC
d8xdAkxS/RTzYE5wCKAHHtmR+PZZ2B4QNjaqq9mMaY8rjjuawrGJwlLAIB0uJ2xT
KxI+4PWIJU9t4DAhgey8o4H6yvYh8ubJ9Nz9M36fCq2g5aqeFZ4NmAjiYmop0SC6
iOWed4k6nfQHXr8i72lyWDNIF4NG6fXTS7eFMZZk6CFOC3OIFx3xrZ6aXFA81F0k
zGyknQ369aJuSkFoIL/ckW15/6QvAwl1V5IwQ8IWFFqmgauGYDgXnM5JgVeWtL7e
pYLHjJGRxTFlTLq4HM/ffixREXp3gQW0K1rAMqsPl3f+mWRPCnVrgyGmTgHBGXwx
zzGZpiscDk2Pf9q5Ter0bb7BABAP0NoY0Gl4ITBkMezriTjbhT8Ep57NEsWhRSao
wztquyGL1vMtyohkvuc2TN7ONI7uGaPy7pZgiefcFaXtzTU23Q7lYzS8tFP6QvqZ
dVYXBO+EVllNpHAyrps+wY+NNk/3f/TvXHN6OJ2Zyq1Lia9agDM9U71W4aPnNxFn
g6wDEFAwf48eRS+YaD5ZSPgFqEqYWrBjr2EPrHYt0IdJgbqJdpUW3Ll1pJInKTyY
VP/v6/+imJaOhQDRXFJFPu8/Pwvf77LEKt2C09Clr1SxceEuSwzufNIHAAi31NIP
k7PKdXC2+rVNhJlygj5SnwTnp9yfYOz4G4vkMf6QDUo9qWxlWCrTa3fh+UHs2UeQ
JH7sF1seqR933PjbuNBRUgBE6R2TzDTrKwL9HN1TlMTUSmRsZo3BoWw1WsflW8iY
nNL0uMwJS89+4jtdLaENfY1cW3Hi8S7a5njRINuyLR9KU3sAHsJTBpbuATfD+dII
7KPl0yTbIOrCamJ4LtFtTk2eFzTViRThd5C1X0nMDAIz9D7ElTvxK1C/dUlNXgMy
NhQ0XhL8IxGe7Gl4tagTTMDDtK99Zm63qGckgKSTNbUyTAdWgmsG6Bpk12pA8hDm
+pYtjRQbTfOkGgrsOHK6ZdUXqsuloasDAqm6rCLnTZdHKsS19FoFOOF+YF1pjjYr
S2yi/HDBywpsl4bBhDuAl2MTkwk0aM1UCgXNwbm2Pmwyf38MJX1Rr6Ow7Z+2R99O
cZCB6gBayxfwm/WrM9Z+FBKpm44QR47oqzm9eQ5NVmKKDNBe6CC52eFQNKffgHQ8
1Fp11MEoad8a/hxfrwwnev/KB4shWhEA7dcbrN/fVpzSbOPA3jOMLGZ+3siJZrrB
CkW8O142dlBBDtCU0OGGJK0AGHN+Y2gCmP6AudD2XvNs9W7f7h3skEyz+ucc7HA6
+7ORTbUjfWJ1QtEdB8QNO1ulE4vgX9Sn7ku91XRcVae96g8t3fffcnvMBUCGT/eO
XbUgntpR8667Qm+cT7N69VE4vaSJ6JKy7MQypLJ6zv+UB8BAE/JIEAGrBCT635cQ
DehnbDTm82Bx7aaLROGOdjqmyLAkhZvTWDFgXm+rTU7lvIjifuvK1nZ/JyCscQKW
eM4LG0iDnElfBmFBJybwDZB8E0PHLFy97Y/SSDisB2Owe3qgEX5Nw5gCiZl7jQ9O
8M6mz2yOlL7S0qjvXrC3mE5DNy+cgKrh2oPUjdVi6JX1sGJ46egeL08o8uVYNcIN
bOVUOQBGwDsdv8axH0gJSd1gcsYbN++2lwuiBZVZ0SWJ9TcD7tf9p9y/ZC3vHSZ3
mAYSyQz0BZqz19IEjkd2oDt8Q2G3n5A9i1cUioke3I/WNNzQ4h38blxUzXdn9Jdp
1frBjZFOtYi1VqHt/lY4e9OUBfsNfbreV+9iKfEmGIGWzs7Pchg7DTT9Jyy353Hx
tmA04SldyMqsNiR0qk3bC3ZHQL/OT7oFYGf+irj3ulEEv+U4/m1ucYKltxNPohX4
3U/O7Oh6pMETDlGMWuOQZxAk6anAThYZgjkRgu2pQfu86x4nldGBlQRZ+GUXUvqI
RQENP2Yh7J/0qmtg+YCaCcKgkpES1d30boiZn0QJ3n4l6CHSygomyf4yjON4WDRK
w1DJz5APREyQhBDTD4/u7vHHSnCGxBRJemdofE1yli33unFcB5aseH7SQnjmfzCo

//pragma protect end_data_block
//pragma protect digest_block
ZZj2v9L4YV1aVFINFileW1u4P5Q=
//pragma protect end_digest_block
//pragma protect end_protected
