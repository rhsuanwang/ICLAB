`ifdef RTL
`define CYCLE_TIME 15
`endif

`ifdef GATE
`define CYCLE_TIME 14
`endif

`define same_id_period 2
`define d_SEED 125
`define d_patnum 50000

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
UBWT9o7U5TlCEcCc+gb8FTDUEWwFVvAR21EJYBWdBRPar6aPF5bHHXpSqSRkeyPX
t2v/B2zXDNi+e0MUC4fFKtrKUX2D4nYoZysSJbOxEr0L0sszliap2hDs5KKhwBAC
B2o7asBVcs7QGQtQmY0Ugk1EIKH1FmiyzxgdZrEQhWn8CDXuPOsJZA==
//pragma protect end_key_block
//pragma protect digest_block
CRmVauijp1nGJ2vH7b5tV+O6zaw=
//pragma protect end_digest_block
//pragma protect data_block
7WL/eJDX9gUYUczKe0thauFgw+RDjTFudbtH6SYBsCyMirEhFl59vL+rD4RYaGRt
66W2XXDe4+JhI5zQPSEkm/Eztc04I/+Io6/0pCfN9JTV1WfXv9Q03jJdPolRmF2X
IGNtbGA0a8VQw4QfQI/2dQr/t9SrXvFO1q8r2Xw4w74+v65/swiHtY4bZiTW4i/Q
byfpRrY82Vuqc+nS+vzG6lv/er/DVP/CyFrNjOZdMigYcbcKGVrb8e3GlSpvcrGl
0LMBobV/hKsQ+FEMRX+9lE6IrA5ZU/wBUNZUvf2+hwnv0+EqY1RhwTYdmfcJmMjO
4il/16ZIYsr/xnL1r2WZxmpvqjIwyRF4Gf5oSWNLFvSilo1snEs3zYBL5PeJZP8o
Z/9+rJugCtCiCHvlbb2AwmfONe4XzRSbj1jBBkJ2PqvbdVsikJNEmHcPxkUPjkcg
CTJYK7mCD1LaobLm0H4dVYdqRPrT4WncnYafnp9GBlNN04gjVbEBYMZfxbSIAuOM
SoCsLx3JCUlGPus2yr+3eBsvAsJn225Pui6h6d2HcPnu9nNhdikvmeGeUvZdJQpb
E0bstZRYJu3pe+I4BWnWdDpUjkbn2rasY5YI0ct073Ix4isc4OfSHvHic6XxhG6R
iTpsFCq46dxa4dpPMUOPJIfTCtV4/ZlreVpficJzsGIY9ZhfrBPDXlHB/XMWhz8b
Og/OG4LWRQzw5RjrV7jjs1Cz16pMrQh/1I/1KM8vwCQAlJ2Sdaml858eJHy2oxk1
KzSLGy4v0c/ObFbSlFfSiABVb06B10SwC1gDby8BGixStFmzU0W63tj2rvVe9zee
PZsl9DgM2IcgJ2YETtUOeuIQckQV/7yVfg9hLMbzGtFIcZ1O66cYEzKua+RGj+08
gZsR3Aq+bqJPb5yP5FewmNjsRzEMZC/cORi2y2m27RzogmVWM91xMkjmjp5posuh
kVpgXIw7gdRJUMsHKUCdnEDE9HfOmA2hStENSPtQmH8m+vssn5qPxISAE8TEyV7r
yc1LayLirdHdSNUsPmyIefbk+ssYBAcqr8PmmUTR6HdwwcV0zrhYuk+txdJCex1W
wM4sPHn7rHIJTzflXS1m5Sa7uAFnn/nH9BplVLwDftt5F8WwKRPaa8J9/ZgfTfCG
jz3G+k1aWhqI+5H/yRrW03gg48lWzgAKTbl8t5eOwLSzGCKSgj9Fbe9J+/Q1NQc8
y7Ta7c+HdjmmaDDyFFySxUd6BhOaILZAdSAYrL+cS3GUykJJklk5Ibn1SH0l8k/X
utvvya2OLUrizBT9yOznZXlu5wc4ccEW8rqeQi42k22za8pYEyRPc8IG3dDrAMlT
G/qdQ+N8Qw0zn1SVmu112qkLblIQdEjdpfsZWzSvB6xtgN2GKIdH0PVLszheb53/
TbgIJZcl5//VZt9yKjUcXKkNbKhn/qumTyZAqXJdeB+MS8I+bu0cVgRt/LfwYExG
CxuJ2pLhtZLCJueoC2dS2em5Zzp+X51DdM2r9txP5GfKw29FMWpD+FYfcsUFz6pA
0yXbUw6qb4kuGFET1MXDFmXBDSsu7lfKkYSI9sGoTTUatHrrQ9XJb9sug703zxqX
xOo2uGjelaLLGloQtI1fJUSZGvKghuQnCMwocmr9dX0ZtsVTPPerLujTAQiMY54h
whFVEbGsbWmhcnNJF6XACjDsOjz03+IPLkR8xAcnHQkYX+fm0sbDWtNEH7KRdxvZ
dx2gSC0uWK4QhJX+IDL7YADFViBRieemducPXtcJzpVyM91knt/xh+/s051s9qwW
59NEMyfZmDgtTqK6XYpyjwNCEya7RV/anE/wzPlRgOJYGGScPD7XerY02sIltLCE
q5nZMr1xPBH4/KZ2scRU5pKbLy6bFx94VWcF5PC7/kx8RWnrtTffmZJXpH7rd0Pg
g/AKu+OFcvyxOB7nnl5dLUcgcSP0TG7we952ZzBfg9HkI3Kj2cWr4s3bw6SLIiF/
5s1VbsvUQ3aQ/CLPbUjH9xsKw3dC2T6vj4HLNQ0d3PSPfMm0tIS4Rx9cPwsW+1K0
PSxTvMSA7+1KDDCZQe/vYfWL5qCxHduZP+YNjgzT1TooI6jk7Ji6xyumKZARZtfR
BB2RKaHOetjjEVVnOFdBQAmqWz7nODB2URHFUOcNuFUS8Jz67g4ssbaJBLUtAi3R
r053yuT0M/cQpVgUjo27sxvs9/FakH5TjAWIqb4GxZNFABzENneybiyRSLNLCkYu
CT8607x5OPjTZQgc8m90nqvAzo6cM22IfRUMOcD3WTXMOHpbxBa2C3WdyAfMQ1kE
DlWCaua97/OaryCa17pOLUFYFmRExpbvF5uUlsExTM/2Ro673z6RdtUjK4hUYBZc
nL61LO3B8r2LbzT+GgHiMbqORDEFe7LBiYgURJZr36Ay6vB6CKq4ZsVmIyxJztYK
e3yaxiv7RJ+tf9zRbPjliQiUD1Y8Vp8K/Nvg7EEOrmb3LcwY+UuISqaT1NZdIJKh
8JGRJBYoF3JRUJ1pNOKPE1qnHE1ypG9GeHceQtcmWrFeQdp4ILpyvQdCVLYQ67jR
pPyNLOEJoedXsYOZOdSBHVpoZy6Nedwh/PnDkf0oQ/RfIoFE6Ia0zm77oLFaK8HZ
xMM5d+Q//65YGlwJPH36RUsuJGg4sy2Q3QXP7CzS5NybyBxe8jfhuXF7RbEL6jIY
/JQ2s4mcKP3qRv2a0i4WsXCkuacFxA/AbKegE0grA6tlrUePpHG/MVwFna0VwLTA
f5Ni+yBl2QjaX/Lb4RWQz4O4nq4sms774+FOI9jmYwf7CpavGBfZ3jyH9n/HPx6A
BrCdpeYa15cal2Eigwgrcbxx9W1p5neQIMsMYltfc6OllYyrt20CH8N/qYSgVjAk
iM6U+noRLhezp4QvLtQs/gwXeC8Jpkcr5cqZbA9V+tGsUVy37FScZW9v+oJ19lM7
tIscHyK12omIIu0FnqbUFDIz19bYgqaMJEEdQlPE55A//m5+KT8oaT6TO/8ketRT
kCxCzh34ze4efMue3RKWcesuuQlvNnzoKW4dwpbL6jKmDeSOuT3/EFREixCL1kUW
KdAKMmZteszM4qS888pgAQOoSk7iVJy2p2skpq/wCK2/kLbQVtf2O68y3ds/rsPi
Wej2dec9LBm2nIpALANDfrnfwYB+Ame9fyeqPwXepihnDvUiE+5Z/WrFodbQFJdW
wcVeMGDAqncKORLdEpf22UXycO52CiCN1hGq6RE07BWEbtbGIH8U/BEn0oI1fG0e
2PQR4dJl3fx69jmOT7JhY+9ONMPBshilv7UM+Dn2Tb8DHjwypB2uKLlwfWerI5mO
mJoElvDWFDPZygPs/FOUuMWy36tcSTlWGC/SESQFjwDAfFa+tkfnsnPkxanUShbT
vo7DgOfDSuWcuFU1XDFWpkw/tzawsfBuf5veaTbTGTJRXraqZgtx9CaliXWOJugW
OtTIb3CayQEI1AJD6JxKZtyMBSE487+zDJ9Egh+EAYw6w8itfjLqVSTWesTQImlw
wmHFLiz8CVGvsab7lAx1pwzkFwk41ycDM1BtyR1OunqTTAvpk93zVDzMxV/OjLHg
oTmpj+sU6zdfYeFSamJvy+xp3Ze1Ynob/24PR2tsidBGh+eWikHQOXYXFdlXS8sz
sgpnkPywiw18T1HHXR6NGWkHBckQRBGOMqVhP0vMljFzg8+2zqA42o9FYmV014UT
dBC0HJh6S0hoWQE8XCFJh4O6BleaZcua4i5XQFnF/+trqR0aM+l5xR0zPuX5UlAU
I74GU6dsn8DGMmJSKHxrzBUaNcU09ERC6B+ioKGzP+gdFLMdzKIZ2LYm0icUyYe9
2OtfcZsRkxegkw5bHjZH/1ZqMhlutX5a8eLe0kqVgnrsET60aUtjRX1L45/H1Z6z
Oo4Fy803qI90A6vTveAXqz17sF4XK6PY1/yOhsFJtbIsYwfDIBBVxWhtisl329ot
isaP+SIZrkb7JR1vwviszxIVIBmv5qQgYv3nCUlRpYxmqsF3E7rl+xGSSRuB5ir2
Ou/ehAeZy2aGLjoQE2N4Unm4msGkqZi2NIheiYl9DNGe1uNHUcJkq3qdBnralmOq
lIsqsRU64JioEgyZbA1n2Di55MKmvEFekdsToeeZCYDlwf+3w0GXB/CUbSfJgZyF
KlmBS3ssV+D+YyMm0qpcJsDaWtXBpKpUaDoD4AomLo6kQXn1p+dCyRGt92oibgQU
65hkf7c6htXA6PJ1VJ1D9+bNMBW/YiGY2G2iOsWa04YwsOHtccppynf0+fug4zQ/
yAeTS5Asr5ItN1qYQgM4qL1kDDwuBE9kaXIlDX+729SRzShOJZTtTH4ZzZk4nX1R
JCTppGXRBMS2MUupTm4czudvGNPsdLX9BlpkIP9tyKlUB3c+LOlhrnwELCC/yN6K
79+Y3kPMasGITO7HAooyVvxeSPsq360BxFmsOdt8CyCn+tzxJz1tKrnEMGOiKmg0
8NwGcX4Gzg2Vqpjpi38o2gPZYD5RLCM80EHgnterqDD2do2zjCcyfuHNWRC4h/9f
WKHPICaB/ZABo1FLdQmF/qsizDqpSNUuFvdOINiYn85LtcyY5Ts1eVoOvfcYVWfM
V/oC9xl6YUBS52rzTqAVbQll4sUKIn54xlhZ77o6RG2wBTVHkqkaLBhmQQjAcpeR
1v7Yd9OJdfSNEcqO3vOCnx/qLu6Yl2VFBAWg8YqWLX9cY0tTkoJSupnrMe80SBHp
AN/6wVpTemQ8DXVMgRLDpwRpLWbYeqMzSHevHScIqzBxS7x2J3TYlZoJGWZL979Q
xK8GUhwsGRlScrB39Pj2KlofBU4oz4ENI7ZZF5lOtY7w2Bnto1ttikaq9ZKDQXM+
T+KEF7bSFHGQ4BJVYA1ggbLNKdsEfl6iDvLcYX3vaibSLxRtJN2ex+pFJKciFWLe
gK5uYJwdU4oRzgCCGgiWFf8Lrxn75siWIBZAjBvqAN0QF3SLQiw2Qty5wwmxJjqc
ajiJf3Zx3YhZ535lRSRiiRxWXeb27B/iepT2OIVDJscUSKqha24oYvbCUnMborYQ
8rMYlNcSp6PeBGdzswFdrs64wxYkCjiM6LGDp1p2hxwyJoLWT1mb17IwQHTHVw7O
evezy4Z/9DTk8tqyvaphJ9SvYcuXihrAIK9efYFvjEvKmVGqNjLOhVI/SpZKCZrC
nNyXoFuI9H/Ne7XesrOBN738LCXfXkW6GOxl+9andphJfk+/eR5QYUUoe85JyisJ
i4X2Ac1FPmwjoRqlste/QyETUUQpGYR10EKsG8AoKM2Z9KWJOCoYyKPOg4r33+tW
jVWl5t2qR47Er2enHlC+KuVoo63BuD8VEIGnukadbGfEDlDmPGgOawqMofjDzKXA
KyKIWanKF+VRhrg0YZX6KbfX5AAGrdQoUGDy4jSkiaei/p89tgDeCZNTkYT/rd+2
fU0/AknSJw2C4W3vJHySrTq5NW+XGqBkn26TGP9hYKL0Yg1whZaMOTqVQlky8L6y
iPF0rdy/J7tR1XWyvifA7hTWCGtUlv8H+ZpuXcFZ+CTKWql4MwZhW5SiE1fexS0I
9K+T7VfQOsYbiAZ1RJvcxfTEkGUqMIea24yv1z9E8NcbD4BUL2qAHX1bYQKzT+bu
FM82GPWhVOroEtJot0zz9efrUpaI+2Oldpuu4mQxLoeUTUTJ+rmUhcB0Hu4XZuZn
bh27w32j7FyGa81NWgPVJaHOdU/M/JkYxWfgxQTGQyjq/zQ/hELm9za7HzhOG10Q
mw5ecW0QobtComO2KbWa/vxt0sOfllOYpJaWhvZHmbGD6m17O9c0FnlUJmRDc9+8
gencnRDYAkmXN08U6umQ5k9HovFVuoFgZbzXE2sDjtTssOUoGoS2ll7zS2hX1iyr
3hiibGM1OdAWDJVk9w13ihvs147cXOxQ15rDGsIU4U3uRKjPAXNnm8o16BN+JkWm
apZbBneoDvjqaeMuJFRbX86DgLlDH/JCyatWpX81QyJJwHMkEuYHPYR25mjDIW9K
LVXnCW0Py5OLut7+l0as+mVfkTQnOgZAXoJ+rlPPIuEXGgpKmJ2n+HMnFjbLFG4w
oGDAH9bJudGm/aNPEWQyY5s7SuNem7G/A7w75Vnm7+ESb2kXYCLui///hnrJhJuK
bVB7rXFTNNMjjn356GXNgx7Xj+wiQ99RGotJJ2TGsEpXz1z8pc0qZegQm350vgnx
dsWSiJbij31vIjjEOBiKQbh582+ppw4OCtHp/hKASjW0Ko+b429oVRKG2nF0hd9I
wz8QZj/a0zzySLT11f86/sdtuztjtVJMvpjrxvoEPJcaXbcH7I2XXjZiS99CjUTk
Yr0Uav1N2MG3l0gwk1C+NnU2tIAoUlCivtJqcJvhaUSI0hfbzqn6HUojBmTVeX0f
nopFyHT2maB7tSpm90IVsAG5cjxKN2NGz4sRTAB8lsUcOAeZygnZgRRj8qmRNdsd
fNe6dzQtdONFOSQsRDVGWnIQ4FKpMiZL/hF7kpQfERhnp856OBQA2UlH7+LNCB1E
1L2/yyU0cGBsac9ZJCuTF2vtdl1jutCxPJ36xJMQ9tW0VPXdSz3CeBtKd9LvfrXK
bLbLf9brl4dhupgQB4EVW1AH4RWyQ5OYQ4VCFIBrP30DNBdDElBV/hr5k6Otikiv
keM+38fk9NRsJcVAfkgmbdkXq0K+0FIJ834dGeH9ipjGbrbt64E0p16UWFeLps7Q
8qS+YvGvO11EECoIvDFGtAPliNQteDN4KDRRpYOXYU4IuqmMmSe3yDnC8xPQgfQ4
xH8Q/2wNiuZ4K9N3CwQ+/ikxfkqSf1K7ZmMpj3gaMALJIPFeBQTOAILPMc/PcqTh
Fn9YuJM7NkDwbi0TVt2xzV9dnKiXjI8ZmLoEg3dasYiyXo5zUw2Qfd/JHv9wE/7f
zdrk6LWToYp1QApkEpU3+w/XJwhWjcyH3wJBnqgrM+CSij5XP1LfTMcxx1vhTyuL
4yVie5xrfmZlchqjKzKKLeziX2c1ehkmzXKBWmi3PXHoy8WP7jdTlHWoNfC4YBZL
TBrI273awgVhIMDFrTB7LMPwGor5kxAoh2VMMzI8gFWkmmp7YztQGZHm6hRISorq
L4H6z8bS+yNIHxf1JXBCgnnVpSxsYj9UhYDP3lnBYyU6ad9G0TcOt+i6YE5fxUUN
SVuEf4WJA5vP9YirlYtKV/lCepUy+YcgfhRijwMjGPkY+WSOrYZ2aVxnFn3oulel
hlP+xOriafZF1tNO+9NQ5gn5JZLe+lWCH6trz/QbJjF960U3f99qLdm/68lyo2wW
qcoLo/OppBbtRNR3OjvfvfnRGMn13ZDnAxN9BbqKJpHaAZ6AvPANbjN1H56mP/b5
Q1xwi8NrN9TrvRfPk3zel5jXQrOT7HVKxZX3nLcwzbyFwAIY7l4NwzrWFPC5snLu
k9sBUqXBDMxJV3fBOiSRZZDFjjH1L0zFlQ7co0M/v+aikZGNnStoCC8UjpxbpEzq
JM8/exuQcSwKiaXItI3XkAZHKfSYmMboPHU7gS0OEjpHReJU8qryF6BUs6HeaTn6
Q++hTA+fvWnFnTc1peLRoYTGwSwoD0dp4p4ZKEl2sushOrneig8bVntk6imRJ53a
XO5BeCDP7W09+rwHpv90AFGCpiDAVznAh1YwoKD/tsxnbCcs89tFicRQwUGX1xxm
nP+cruHjZTS+whPz0xp3iC3cEWaNFNJYOiUH56srbXu9Z7t45KT2X8kEo+KDqFK/
3Us8cZSzaFphAJAItWMmk+0QzHQYxI6g9AOVc/6N1+0X1jMtO5xQsdV6mYqHLBUZ
RWUgYlE7f/aa/yJyTrkSaFaNghiUDqio4ZtCplkqRlWjYSfXnf/akKYGZ9MJLDNS
cqP9LRL+fXepTUTVuhUQKLu0a2GDfZfNLsHh82IVGQNvwa6e2uPTlY5xPLpHW1Zb
WU9qPKbep/BtKrgbVHBYDPYEXizHVWw871sMU7slp6DC3DEPX9Ojxh8VCoNpsSjg
eiI1vw0hVcfOarcGAw4rTW/pGPiLs+iMBAq7MqeJjXaruhh2IMXfdOXq9XfIXE+I
+7SbIsTI0UeHHjQAy7TJAnGsUhamGgipBszoEcPC7rr5Cl2S+9NB6r6quBISN6vU
Lwej/tvXTZ735pWRyXYl4TRk1obZ6Fyp2fz4KNwjxmRW5gwB06rxV+Ey+Cax0K1w
jgMl+6yVFBAPmkCxgIe+zrasnI2fsgKdEhqSzRlYAYzvzxRxQ1muv+oVw4yaCykN
Z5Ia9m4qBlbrKmwJZx1SFYRVpCCM/KGQaBz75jGi5sjeBH5hh9DLMBo5IpRHoPN6
JutssfFPbrkAdjX30cC/kAS1N906+3f6kFZlga6BkVdvAnbj9smZx5yIxwZrXjFm
JtpG6p0rksy9+oXbAu/ygo/mB2Tk4ScniEb/e1k9+bCBEmaau4nud0nErnXWQC6+
B/T69ryEyXKCjjmGBvHow2uwA+76Zx3v9PIdNkgTeghxr5ok8xsAD+DqR0ET3iai
eqnNAM0mqdvCKIjnOB0rCV9Dq2jUYgznpfLT0MzHfj1ALP4X4ZKBnzlBr9jXwbd2
sGdl419g2Auuz2TXq0WBqFJOcAVMCmg3JhhloVx27Ik3+irKEVJjVxaXSzGujPsh
c72+P+6lRjljWFaM/fJZMnh0sJDFcFlOlN+PLnZbuSigkKakHSpW+0gNRnk2P73P
UYqJSWgAy6cIvOeynHy0thvJNMvduNMy1likY/gMU9pnRH8yN2gH4ZnYM0oc81oy
m1fA2VnNoZHUjGfcjcRjB9V+zyGporRDJclSMDic2pOcW0OJFNNVDRX9dwexO3op
SKtF9ehGfYa91cVMscAOGDGyyC4bzzRllID/7eNEQAB7pI27SSN06Jj2zUUiaHus
J7lNJanjWz6H/X8i95AHSEjCkWBIPqSM+dPb3wJztvdZlf0dGyTltnsxOXWNMEJu
8VrJTFHi/wHCDYhFnwr2SSE9LsIFqr4mcxcDKJMxF9OQ2YEzoMXN4krXikvBaZDe
kCv0pcqaywRkbLg5zBZHsILWgKuVydgeD2Sj6/fIwkpPrlWrgT9t1lBJYnlTU+W3
mgWG35W0TshU+F11H+JYcmjJJHPA94amUjhTgqk7aB8lh6dr2KU6s2+KP52YXo5H
sIiZNcPzegNknCtJ4fHXbIELXxaUR1NOMYJb8gh931pVygn5CG1804l+SBhiJGXO
c8azP1/rWqFec28QpedAAn0EfRPnjpi1oE3smhtzoE+W17JW9fGL24dO8FW/rljx
YedAzucggqjKuuZEKEBFahc5pn5fb82ggzXxfp48JSqqE3Z+iZT2JlKxsArWo1LJ
JqYT/Z7OHePua8cupq4ejq+92myYbgkZgIPnnoWW6x7sz/9HEDfy2CuHnAwTl4rr
PU57aV51wa74mDIlYzOMMK0w8SXl0yAyzFEpLPf1M1KVNKYW9P/SmiTVL+h/GZPW
H48Ts6qtz4KOMgtxUBoTkk3KNx7zCXKVKpqpk2YBwVZFaG16HnPiFJ2lz/X0+pvt
yOJ4geThlnrT4BQUThbd68xGDppINRBbRKp4z3AghWLAaZpVwIRAfSVfmJOow8hF
2wdXaEkHdC/ggyaD5gV+sPapYzJhRyZBrGDg7Iq8B7aTAOc7kf+xBGAEbZf5MbcI
Evycn1M/QbInfFMhMtDmCrU8M/2SBYbl0xTA8yFaxBtIPrV2ww47SaldZrQg8bDb
NBh4BRdKyD2vYjwSetTodnmxkNIRtZYW8eFugmxD5D5+QB2GRJAWoMHtfWXrXcxF
iaB8brmA/eMGKBlkC7cpMkElwJ2yh2/hPINlXUIqI5hzONTSDgS8y02v74A0ELFf
jSwwxUpC/gZBYKT17xeY8yMAS3vbjx/OzCAls1QnzIgJyYu1lTGYNbaalPz1vymt
QFjrAbNGm1DXJyDjG5RGP3WImdUCtZJBH3A07504wcvGcj1WRYwLtyJwDAmr5Sn/
hdX4U59q8kiIp7jArJEBLF2UmsGInnDnWhKr7ihZS7cA7KhP0LPfzTJbSIrVHWON
79ZBzde0XY+6H8awdveUGo8+xk7gVyOs9KSZiknIVmIlG8cSystPMiussnRv/lPD
jol7HAv3nLoUvZdJqpRS9q6RZm3CAV/DeckvhF0T83vdgio69vP6+3tuHl9xHH9x
w0frnbrglCNXRzVDYQmAswKKOQzIhe/J9mU60LMFnG8I4NyOqJjnhaspy7EvvzLL
E6lyyw6ImOeid30ToLzjEB/H0W9R5L9yYo7arG7Q6W9otnGoZBtxHJlyCQpHAeA2
hFdRHIPHImk6bcPtjpvs5t19bbl6bsdKP1r4YPonu/VY0rmHS6nwFA+qSC0/7lWS
qagDj9DwRKh1De0k4bs0z0jxgk7YYVnIrftX2zvj1n+90vcrdkpjlamg2cKL7HSa
Mo0uKoEU/N37y0ANWKaFVZMS+USAmBAj1m3R8uMf4fVYbwsYYg3E27r0BObkIkk7
Z2p0X1Kgg/yzQuaEFLh7/rJRaIB9wbu5Sk96BUQH/iBvj9Me6ThKPgVy9gFRrHcA
eDOTSiTRg0y4vzcjcT0Weeq3yYddtFzuUqw5rxthJ0vYVPb3VrX97OIpoZPFdoCK
CNLeOSrgO8OQfTsaulYy5ZjHez/RZSt9iH57DNcXScxa/XDg2jUB5aiBEaEwJvnc
YWi+7lEyhZaPcFFwgfIkhSLpr3ORT9L9hGsIiF9a1k+RkEXiAAM/nh4iY8kwz0tA
p+EdytJxt1s3KOTm+/6ov/rj8ZoxzWOpMA/zogsxZAruqiQG/pZcThIOG/78JtOv
iWXiWoANpUTc3S8oltVFFQAgN4Dswa8HZvG2qnIAMHZFu1OV/VsV17psH7hCEM8h
Yv0TATyAJ7phIx7H3JsFy19fNCenbdUmM8wjMeCWWb5iEuXAS/FUXyObhLqKvlc0
UD6r+xs9cM8gduzpo+H/T7FNJH7lxe0yNT0xrb/im9TSH6LC9ipxmyJZxXqtQh69
dBx1oUZguZ/W54/Pxxj4UTHMhqSQAZgiWiAjz9o+zoLjITfprS8xmHgZBQPUsfbW
6owJZuYmSqq4wyzBdR45dtLmuHo3lcs3aC192aWmclPABh7GaOQkeHzvFVa3c/UY
AJ8lruJWn6yVkWUBwh56tbWm2A8L8GHZqK/Yw9vtykdtd8X0lK+N/iNJBxVKKebs
PQ4nsImAk3D6tW92nuJI7TwCs0igj71MclK4S+1mNQxqCfRhRwfFOohH8GR1m7Lp
bzXEFeCRsQVo2MGoY9v3kcj/ZnCmEeQCfIL+OZdcJL3GSqR7DwUyfzFcUk4gA2bZ
gR+cp0i9J1U6c9E71KBSixKzRnXLerGoRypkc3ITUzy3YJAGFeaMs+aAxFIvBbbd
nMS2AuCv0xhGaKHlQ+LRzUAXnmQzSp7pg40PXyjb9VsxmeuwttnZ1G3ovF9c/byB
tmqtdaY9ojFLfXbo0Cqhfl8By0HXD5KXCFbWrbXN4x/gJi4kbFIKZADmoTN+lK+b
X55Ic7023NTNXBP6WPI7hZIJRQkueiAzkc1ucY6Ef9PvgHVxPIg3hgwFwxwD7iNl
qUFADDg5JLug/J+mw9Orybdg/GVlnf2RVd+sCFQLy671S1AkvLjh+7s+24I6uPki
OqQqvQkGxdMRh715ANsS5ad6Sv5IEZPUa2zBdu2n+u0eBFqsF+QnAFWbo7N0cXf4
cdJY1lkKCi+Bk3GD6G4MPbp83ytb3uHaLqUa69s1Ht80QRvJTUYA4nDCPe9y+TlR
9CPBiaZI3bGyjYBcUkig6PjGXSY0woAlqY9rEPQPIDwT8I7zMstox4qBlEDr0Esa
lodLUx2wAbj/jcuwBn5skWTkcY5uXZnnEUS8rkvRxt8/Llzb5GeYdywQPZSMO9g4
VIZjd5LhjvYr1/BUyK+mbFlMZx+cuAkjgHvOL7cQ4L0+CaSzLv9JfXlpQNVOHJwq
ADJgiJG/fmYmyEGZUrNvzp5FpgzQrL0awXweWPC627huA8ZzmrDCpLoTisO2PRSi
9IjZsW3gNUz6En5DYoArv90aRhw9DHmQa5qfv/1gdks+J1TF14ThD+EQYHp+Dr7C
Qw8M6zweBkk8onCdPdx1dpQBjdx+Mpuwgk7CnxN2fbNrbn9ECrAb8SREHW8EJnpc
OV6t98Ypu7sJpXLHuxlrf6VCaPLyZBzzX+y+9rdy09qvNKCvy8RifI7sJaqelJ+v
UhFzeP7rsETb56a0fwhoPuWbfknv847A20Zq3Piz8SqeTpWxP05nwz6AWzylI7zv
LJ1Ich1G8j5GUX+/d498QsV8TZD6pKJPOvaqQ72KwY+RHC3A12ST7LzSqBl6qcwI
WCEXRDsAVUUXnuRlNlMYntOxjUcaaM4ESAPk3VTx76ZENZHFcT2MTQJc1HUwiD2/
9MbDdSgeCPAgVX7cckypWBv2nwTzoybu/KM9yIHIp3woU4h4h/xPVsh69iHufud7
pkxTrur3Y11+cW5XoTbcPSJiva/FCE/kJjbBvCb9N2vjryxDhkvXl6Ty48tCy5mN
X+g62e8gCaYW4Axbf51kqVUbVGJaLh2NmzilS3g9DOCOPlOXe4qsH4Mj2RbdIczh
Rns1z1JSqi9Ci9sxCctghRs13YFnnL54waN/Nc1DB4l5wKtMsHvlLtut3HKRkevZ
vMPYz0aPn5Tt4RFLxSfDbhrkpqd6VMzcveLETSv0YggO7TcIShtWG//jDxACFwtZ
vNowsS0Yxe70Vrk4igpMx6/nYHXIU3J6J97rSH41kyfPWxW4mZ0RcN3K1EsQ3FyT
tICts3n6mdt7sfA6ShanSFsMsNNHrXmobn2Ra9X+aBVq41TbCaRxRmUZwJs4c1W8
/Aus+7kipYQysuYC59ZwaXhkXS5XNFrUuyF2qNkgZ+7xdXg1EFhu/6uLtCFE5gga
FZo8mtKlvCls18Quj2gbBlpkelcdp/ceApgOoKX7BoB59t3LROvyWqMPLOC2KTxo
oulIX0F5f+9skFwXbk8qPsYD11IeEYitjB+H+RCMIsI5ks5mCWESL4Ro4eItECjy
O2XzUYubpqpUStRQm/1WeZ0ro3uGAT+B+f4jHo5b88zRtPjhmi+P8y6PXZjZOLje
/EShnBJRORXMg7ZpMEWqtOvB+QZfHUW7c6RKewtXSfnX5A5gP7Vj3XcoffmfsHt3
xvC8/XOWSqFqlMhIp7Biov1QUcltymDDiUugWIU1Zqu26gYYUrA90RK/+H/WtJVT
qORG+S8OaYU9jH6udMOOpyaTU+BgV4nf3fq7k7tw5guTAGdSVHTWfpo7DMnzwg3W
P4iC+kjd9K8hpzriU6cMHWP7b8Zg6Gy7npjW5dZQ7ACL9OgjPz4gwcE1o7RXaRMl
KSiP3pKNGZxS528anU4TCj1JJ/Cdrb9X1TrsMry1uFBSiXafspG9K6PXhxIIRub+
JI2zqHv7n5lGkOG2PefZglwkBZ99zX6yZ1olYas9qNI9hw0FnL9Kyp4vf/YYc9sI
2ReGqMiErbQ6cYbajldS6GD/pzQcmKYy/cJZZKa3LfdLTZE3fksJqVYHv7I1+49n
MGd4zmkvcrvCxgI+O2RZbuhVeN+Oqfa/LAYT+/v8YHCxFArnFO0OUT+JaMHQO1YL
MxS0N98NM6XWfJrd2dd1NHBt4lnkfxoQKXy5cHHCdjYAkK4Xk2BmqaJonVY1gN0Z
xdIzlrpf/ng13cXoRRrsUVpLluALXoBVR/fwWZcRMo7LpUAxd1VrdDWByoEp9T2y
tN0kzBH81HZbdgb+KJ77coezC5xhzViJvz3/QO5Cvg1U7zlcly/+ETiJkmfacGeD
tMyYOZCgjYuqo59D7XMkfPL7BlZOhUwuhaoSnE7pGdnkMRIzUb5lO5L9KoqwfEfx
/uaP59IiFpKChJfWZr1JDLAR3Mp+rxbLLdjs1d6cRjabm5hcT8/glrqYzPvAKW27
1PIa1RscpRxCrUmpqqZv7+27TTTumv9frzhL7lv6zwcP9OeJAiGOSP5VDhsoNz5R
CSpCaSAOBYfleiU1bPiXaFAgLOxsNCm7/6Qn5+NAh9kZ6feWjLIXVMhDw8da3cFi
4uwuQyB4yVuxVxitKvfVsUV3/epiLmkUPpUNP0brUgxNvFtTq4TPwrDE+dIfdD9w
6zE5HGPoSqdH+AyZL/xSHZDf2XE0+HUpLUhcgXxDkZrFZJ32nN5hKsEAdFe1YmaX
5pC4mXE9McLKYo/OgwR4g+S4DQ/zXwOACRL0MYTrFcHEM9aMahQ49/J2pQs7PqEL
+urSxqCkm9K2XRudOyqy39Fh7f9SZkwE5wxIeIoFPz3fNLR9OrFs/0Rsd2sqWGaq
enB/KiPwtIxDXku9d05qN2kvblofR4S8QnjynPAAO97d5RfI667z+AzH8oa2EaL4
vWmTYx6bVuNDXmLQ7a6fRlv7qaLajreT2umnMxc7x6LAmYVJY3ThNZwdpDvpZxTW
bHWJL5UxO3UGKMy4grAVwWqq8AClXM2hIwbzORz1HZp5Bbep1h+yhU9Z3GIFEJ9v
kSP8/EUxOOdowTBWoDc8tqopbfQpkT+8TEjK3zr8z2NbF9K9BWoSMwxrvaqqS3Ot
/XVkSHr6RBW1FBuJ7wAEhvLKXAO9w2Nga4rpddATZWY9J/I7/m6cEioGaooRhuO3
qPArEWGiCjWXZUa2XlMN/hhi6U4n1qVMdGB78ooD89B0zXK59p29sr5l1AQasYLH
bSGTRtb9oWcihIt4td/4UCqA7w+t7ge2n4FW9HprbT1AJ9EwnhXvzmG0HhcZfT+0
K940FdzMkqePQ7D35HsXK7/fRRo/MMmvl3c/2ruw/hdQbg6t3mpceFq7wPFfqOji
ypVxA5sEqOo+FIxQc2+auLOF1EFYRuZeqjFBV5y6+CFw8B72wlmH0t+KY3lqP453
GBqGJDUXpUUGJq1ZXKe1NjPzYxNrJIr1inQqK3WyA7ci052fUTEMT4Alv7OOAXsY
k7j8l+celDTxWfjMKXp8YlGsPnrFQPSCV9iGvu1ZnCXBkKrnzccIURsoITjS42fL
l3CzySw3lVvlj8xxpvnrzHEePL3FK+iFKSaEr9lKMUF/v8tC0ykh5zO2AmnK8X+M
egJ6u7eN94qBtoLJMsja5dND3o5XsKMeu1aQv+HWq8US8WHiiNFWro/NvpbVa11j
Tah8WRrfRhfk84O51ggu8u/taVEHEar8G/gjb9C9+FG8HhriuBRrw6TeAR6r9Tyz
SQ5XvseNo9pSG0Sf9h/2DEvw1isMuIAJpQs6c3pPDtDT2BrGSoRqwe54xEk08rod
OvteZ9KdSVOlY9U5VuPmXwKVQlvlgHilNdVPxT5PpGyn/igaPHLMguZ+t30dFcDx
oXe+Q8tfBiKNAd52+FXCzV0eODU3deFSXIeKMoDzzbsmXrZKOaWAU1o7F/Pl85E/
+hPxrsIH1791wm+Fg0nsTJsvkiIdKMFjVVks3WXLjWW19y+Vy14Plhm7vRDQ//7e
qIl41YB5P3yv9s8P2NYGTllyLd7+CXdlqYZQpEqNKqVRX8bYk+Kmv1Fkbpe0093y
4xRvqs9C/28AljGAUXxe9HhanIhgnFz1HuQ9OGseC5mXcJoG18wt4YcV+dBa91iw
Q9UiqkpIiCQc3SrF44vn/wLisN7NYETqix9F3cFylJst1uaGXsqF3dgcTgvXxMDh
JUs+/pf40UegdDYh26yf7iwerfS0n2EswvZfbWBjYe3ukbJ07tVUM1Q3Mps0/2dd
wwVoLrkEg6Rvhnv6QxaBurXP7qs3tbuBoOK3idNRYx07TaBKISmxA4B6AySyZl5g
9sCT//pDVUUUouHHb6ofgLfvydcrX8oYNdKLH2kuUyN6dXH0LSd9QhtNos16dSgD
PCsU96TtgHQJE8hbP8fSTujiMRZFpiLo6NgUa3+aR/icURkgSV3pieVAJwIuPL0M
2AirZsqHcZET9KEOteY3/sftiliL/I3ZJ4ijKOr8w1P78v1we5GOg8Cezdlh94mA
5wwf10Gn9448YbGzewdVN9JmOScNut+yFaOoIAanZjrryJivIVr+u9TKdwq3vp7Z
duQidJzxrsGNSkAZSYc2NvMJFZOnF0YPzk2lkSMV2pH7qDyHvzFpkDMaCTyREwUs
l9WX4xeL5kJGTrShwLET6rDpPox38BFbbg2OBcIwDwIMqmGi31M1+dgRmZRA3o49
23VqOFR55FP8NlsI/ZYM7Zp5HbSr/IiBWauquMf+049KeP+f9lhEnh/A1KV/t0Ql
4hw9Wc9vC6z0gREGJsuwepBXsTjrp7qcIe0wqmL6L9H5SV2vo1T/1RjETrPwqAMF
S6JLYfMom2hhjrjvVfjfgVG1z8fKZO6euIYs+1YxMoBy/ARy4ol69Wo6SUA3gY4U
dYmKeHQWynlhb2XEB9yuU4Ya60E2bNEoJ1emc4jZoKKUefe07WMYHLpi/8MSqguX
4vwBtrmwzDp/i+QDkfcOLaWh4xvt2UU6M+axl3u/0Trgcx+htBT3vvTxywvA9G/4
Z4oKBtV4n02pMN6ogxm0EDVDp9U96wJPg8NyWJrnvF5uuMD39A72pCLJR/7iKrRO
bllAI6jzqOj4+3Q7J8C7dCpKgyN9qsfOtq0BJO8itfD4jtJUn2gGzgeXHhLuN9ru
zLs1XVye1Zoex89s0LkDDf+llfxWj5qNITI7/oAndn3/ckmIiuaAlkVq0+0WLMGW
ELMfEVAxF5E+RQYFeyJckHIZyZY6J4B4G0VwnqHWMqIboU/lDTxPMQfYt5i+lQI+
c4efjN9XS1eaGPOt7p+ATcktPDmvuzj5GDpowGPAKh8MA1+8lb2NjkhkuM9LvOxp
sfwIb4bM5Z57izgTRpjxyz9ZtRuJ3slq5Xgn/8NLIoJvUoBAlZXBq38ubM3uTBUK
oKWOnof/wewSb76HWdzhij9VAlpkRhovZ6fppA/MI9i6KNodK9pG+hdi4w2rapPU
e+QvuefdnM2O5h+Hx24c1gSUK5Gu78T32MgYY/CK+wPG75NEru2PWoaX79vKZVpF
DXvDpASQMmJAQ+42Wt+G3GYHnfTC3NzOvyBJ71JHwibYUyscP2seAk8o+E2J1Vgk
kcZBWRIRM2WaqPxFAqy4+eBQg/vcKi2T4P/LTX6dX4/P9/uqxK389jl/ggZH/RWF
YnUfPEi3Hdox/o/opLl/y2AUXEUXSRVQyZuRWIZOtXOhQuDwapqzTAZ4DstdE6sY
yHNJjUlxxh1xNkmykAAYlb1S9nshdA9+3FmdNiynjjw4Dn3m22YGGzSO0pYWg4BT
QHSkp+q1b68W/rX6opRPyCAyxik3fpLAP2qsSUmzSVgT4qvkG4ykIfQBhpv+yHmE
4sZMDEhb0unpJ4T1YBgN0A8ti/01vMqQCfRGZZE6S3P4rtNShDxxxsm3omekuFOz
GMaD84zlM2i41eojlumpD1GuKZ4Aib3TnrRsdW+cpaRC+MTKUSvO5iwrK+sv0vZ2
2Y+Q8+GKS4OJY/BTshV1q8FisNckLAI8p/jl0oRzFMwc5P2Jro2RxtSRQK4OLnHC
UmQXKWb597AA0xojADiVBwoKCJESM+c8davAwLX1J0levxNxbf/QGK7eSOt2l4lh
+Q3JB6kAjsT1Md1dR4LomRnboommctCn0Xsbla2Fokgid6K5ODiVXjmd75SvSvPY
aOGIV37nwFrz6e1Q6UQ8wLnHi8O3t6ZM/JjJ5zofYmn2Q7v9gW2YxqlVLyi9WVr+
5yhP2drRPIoPpZ20xxbbp1zzGfJDZsFyKFqM6uOoLO/U7i2EmgVSOU8aZwsyhypk
Cu8vmC1CFJb+UJtR/dVoct0z0ant2FUHkTWPeH6nfdAlzRBN5jJ/15kmpMc+DU30
8U6MCOtq8I7LbEHrgf2P8qs9CQ6VP28VvESkBqtyDpQOsVdK9/OsDpgqlF/xaDxN
HggsPx4kq2w8E8VMYLbHw7+DbkelMgURayDycyHE9pJDqv5BbpKSQkDNmzZ9mmka
sCXeiSEqXRly/OZjt2JHoMokf2vAVXJMuXf+6NnNAmkUg3SGXQT6U2uhz1Z/UTJS
7sjkofoGusj3UpiGRC/Qg6BMvHgNj2bfb/r9r9bTNF37l4B4U9SG8NHcycMv8GzU
1wOHCMC/TLzjbkHDZGvtpNTlZtoMaJbD11NBEL7Vd57xwBwBOSOkNwRKYAkk5zQT
eviaNB/e2ZuTlZzFYO445N17hkqbH0q5xBMFfiMpArNOuKNQGcE+lO9YzuH0SvNq
uZSCE9wWVI34XHkUnbazrDqwh6YnHL/I9Tr9VOrF95zsKQmQwl431ZXl1bCFH4Lb
/GIR8UubWsVU2z31AfY0dz2soszWfyVJhEaZxH1efA/1g8UOBxxvTqg7P11DmfIv
VZK3tBB5H/vQ96dTIv5Xt6udrCv67mFxIG2mufMmpXUOE31lb6LnH6BPVBPj2ps3
xcWQmKvVYon7YCpasqxdJSCJngifYhKxlZ4jDpyByjGOV0SrUEYeLxi7GQ8PtsET
BdaLkBU8QTIUjWAwccXEdXuD2nzVLSKDz/mRxnQ9/mY4ZK84i+Pn3O9bX8yF5hs5
Gqlr3nxMSJZnW95XIL9BvvHbwcCKr8z1/xpxfi54uykdE4ZGwpjC3p1KfGJP6v85
XexdekS2uNq6bnK9TKcMqBY/V397h/WGVvaDTFYNSDDLxCScmgjKY//4hTEC0l2B
rfbEaGHpN2loHFbGHBHE+TBJr5u8MuwpfDKYgz38ETdUj1JTFOBWSbOB6saDb45b
ZiCt8Pn5uIUUvlOwrbqOf+pgpX+KlgtLWIsR348+6SzD4a1+/9hDIi7Eh60L9H4B
SqiREwJxbjIihlUfcReis7N8lV/0RY9j0/Na54zRZ6L9Wz8PTdqwYrCXRNiYftkJ
wknUsVFzt2Id3GcmB5sYPHy3wX6DDOiVwm/Orc7v4mOFUJWcqabMvhPMdheuK2xo
nq/m2KfY/fK6FvdtZ/iMo2Y7aow3czk7xfehUP4KSyaVNYsZWHMX1xpYFD2uw8rT
Der1qLKax1cIsB8wiRQ8cjKAhPwchzzPnEmVwMYBdKQujmkubCfyq3WVGZwLmqSh
ipxY1otBFyWIquMe0WEKeEa7ZKGX8XcmJzNWZDWsRZp/AYJ3LiTv5uSWyhxbOYjv
+etzHXHchsGWHXLiLJ8Lp5NvHadcm8v++sMnr5e6ov6FK+IbZAzOuPIXCl2J9fi2
wgYzVEipu747gIJK5QPi62BA9Q0OHZrgCNluS9fAgw2pnOquguM8olalcBf0oTj7
u5zdPKRYdQi4zGB4Iu1St/n3hf6+xNCDBBYdcot4R5tFcSCF4O1AsUzrCD80GjAY
ToyzBxae9Q6NpKzkCUr8q/TZe/z4xNtMOU/s7bRJuhc9kAIKbe6aqbpHof50zJAt
RILrsQb7zPSVy8XYv+hHMdgz7H4PP7G/AIEE3KKsQ667UTuVVqk4DU2HnepOA9uL
hnEtEbEaggcou2+CbjYnW3sPypAFeNJetYksm2sx3V0ky8kFVwS7ESd0fOKE4GXn
yTUcS545VegdsJLNg6NfwFcbgsvRz0lp44gJi9MpLj+TqEl0zx5rXjpdkKwcsfGj
UtZHIBgl8fT8uZv5Yxj7xbs+bWBp3+veoD1cuyIQYmMi9aVRoHg2UG19eFpAG6mw
AYMPsWVle37uQSLAWifA50y9Lh6R7ZGrKjkzRbPaOqNin9E9hc3sZaIH6i0wjGu0
+ArPdrfoLLzl7OxJzY+y1FVKqvPkY2AIsSH1Aacxm7pYBP2FLy0wZZI2mf7NXA6P
lvSeZwLZ0TGeCO0LjVQLIALwTeuSgAhEKfG9RVbM0mSsWCo6YU73XN2l4iI5CnfW
nw2gWsgVrHo6t4kUnbvZCOXsmC6WisGo6xXI/GX7jOHJohrWSJ5USgoZDt0uyRlE
gePlk37KdGz+tOZljC9Aulu2DrtQ2Z5O3ljxBspegbJNhHzQraMhzipzqNayZ++T
Rlj+aIz4OrIBhB1YzhyBZkzXMp7Ki7Lra8iv3lSvKT3k93w6vuJDkZDBAeAXILvp
mnO/DmcdyUYrXJJsSKYruUO1lMoBd8j1eUtm/4x25OhPhyPAPOp1uPfwJMj3DoG+
2DSKCz+kHKmlC0/q+XWDyhv7UoBg+bMaAX927+/BJ1lqLOGxNRTDsFxQKfPmvSTB
+qlgtaLgIsIfa86cnzRtYjR6qCBAFo0N3noH/kktNXuT8xvLtV3PVkBQ0E0YSZPZ
5Qtp2G3bVtF1URsRnslq/tYtkiJXl22uxpm1HyEy3ZF7ZqvEwlGqgu5/8MNDUgOm
/8/v4CQnHrYRG9ODqsqtgSM72KCiQIDgayvcuRe1QOkdtpMki0xJz/aylwXJUf/N
8r740gwEFIDSWK6yqs6iZ1SKVzn+eb1lZ4aqq1pvIw78OCy7GfPq40fQWjXkoT5B
jt3lnAXQcJgRzCGWwMnFwh/8vIujU5BPRMABymKqcUZfZ0CdegX98dRAg95RHtnd
VknqwEtp92YWskZAECMuqdLvT4aa+i1Q8e8LDGz1ijtpL5uQtI+BSrayaZPTzI/u
Pot4fQniT7Zp9NF5eA2v/Pmx8EK8lEZaDaO+Zhi/eoDTz0eS7sq7ZTROvEf4uLQl
cdgk3vZoRuYMisRR+wrx7d0+tCFBYPbNXfruONDr6YhPgiss+dfU2ALhvbR5s/4i
QEKlX+g4m518ZF1hP0BOZeP4/sVRqomzHNCEDjqR+QXQctZPeWpjBukEGoNJFwwq
0g1frk5pp/ne8x8APpeLYdGxsR+XBnfTF5+hsccvW0LRZ7L5VJd1ZUkoZ2t3arlJ
GE/yBZt3twgjGxhXQ6sxq0izCFjncpT50AXQ+AP5oIR97JaMP+y9UVknVvMsWx2f
9BlM1fCo7FDeEe/tfzRBgxSpWy/HfTecGEmARKQpNi9gpJ9bHr56jXaRabWmphds
cVGN2vEQC0QBvODKqrtyEDpy2I3e83dOIOQvUJznvhvzwkHp+nGnIH6MQlZTFIpQ
sbnOEHzgWMyPLBbfjp/vWFiYxaOJQrwDaIm9rC7MqpLTLKy4ajs5YZE1i3RDdX3J
7m1QVQLsPk/VTCA+tfMWohG4K2tG3V4pUG9guMybwTvLhSjdyJh3XMmtgoRMVV/N
7O26XjX133jbKzYkEt9aNBfk7W9qezJ8cXuUpsmIVGS5bYpBbNyKpBDCuVZ+NFf1
ToPI6UWYjdtxSgwFQYjuR+9CegyiOdjoSk/HQGB8bcOtzfd7eKdUcefFJX36W7Th
pmpCBPNKI3mwQ6YJLjjurZrPiXYZIO7QbXVdmZ3wnsj84Lo3p+UckTALOB5W0xw7
dT88NO5LqUjIjKLKPesDLk80v9W5n+wQmzjtgNoyNisbo15A9z42RE9xfwFRow3X
UNMkapvemiI+EIPH2h/JEtZbXg3Wjn/+buyG+hRNiJsEicaQjSiI7ujoELwTWRkc
P8BoqofJqBKj+OFCIGGocdm4x7KrSpLFG5MLwpv3BPDh5oflQpFq/E3yaPc4NCnT
xsWyVwRcLHRnFWMOZ+vXhJ2kCLS/48VLGSG28RykSG9j3WoRXRmg1HwtbmGeTRM4
rE1jZcGEMaw+zZM+VqkgkrqdLBJXHNf6wQWJt5n938rnAZrlI8vUa25faKIBbXXb
drE6gA0ea4ft2+cYHxAEMDh0Skk0oW4c9H/oXmOvsAqULD/8M19OAhtoeozGk6lT
mXptyJPg6dejVTv6qP/4e/QPsAWTg7O7d/y8sGGFlIuV7jql9t5HQOcUj7IX4K89
xPBHI+uSlvfXJEsQ5TRA0zCM5rjfUNQoJuAeMJkvmBm9Vrij+2NkGsjHerH2rr73
xU2zt3THqZSz5mRHw2mwEbiPGiDiT9oIoXQjepRqaOb5l6Gibzc4UOEmUOQyuJSD
3lO3QA0qFzhGrtQAkBnANL33AVfT4GOTDVexyu6XmKkLL+bOa79YoZ52PVY4zDY6
iQPf5spjwkDNuZGlQtSpBorf6T8rv8ruAGudpGNKkKrp32IdBDmHHfk8hwQwuWgm
RIeI9ceZWDdz56FGhqOPMm25Ojw1hRq1YG9OWISgkemiQkJ/+KBvFjKmI49HbDqL
LZq+REvHN+nlXaknmM8BCvobBk0BmNbB6jf/oyKTVk/HFcuuXHaKjCBD6Ru+5KB1
mGt+GZ33CcolKFVw0n0OtsV9iD+6l+9sa4wQ8HIt3h0z5rDe1jd5Ez3/IMRY3Xo/
pP51ZwrCcfOiH88eToEnGjbuXX8jnokUNFuiBw191VAKk7K5H43qjDawhnWFFfH0
9WRF+VS1nt7iB7ZkOu5+wVSGgTTHX+yDh2fRIzmhcBJgVQb7pnXlCN+aC6AsXWfD
0qIYXzk7fmMT5FVw2HBMMmSWmd3rFMmnW3OYCMnVDqSimPZZfBkR7qem/Cwy/GXu
nPe+xd2ORA2PHmBfksj8Ga/8AbvgF6WE3LlhXdl/9XHC+IEGZzeVSWJROnU21v2r
EtwQvNNCvnQUtBcA4QU4yNxrv71Ad4ZRAGTQHv6vcQAVKPgs7bRzyAJsU1nT1Bdg
J8DoHb2TwTH/EvV+y48wZdin6oufUQ3F4BYlGngCv2aiRWkSPGSrc0K2/QCqu+F2
P1OY6n67wAiCc3A4ucIfjscNIPuRxZ6OSrtWP8879NOkRChAycI9U9LlFsQWjzTo
vxeevhfjKLx/BPrYDI5poM7CwgGgIgvv3KOF7Xtb0R1USlMH1XNXR8DTbYPk7DTT
V/zNmWe3t6qoZm5gTQTao4654wIIQ9uI4CtAlT2EzuhkQ7rb7DPpGYMfilO4hGF+
IRE8WLkGJOfq+0+j+VIgnaOuSOmFwnHJM1yEigwfZxCLcB3nw3SZYcbH1JvSB0VC
voVpyg8yj/ioEqO/Dm9hPcsD1MWNZRbN6g1XNpYM/3dfwrx7ZFINBRdDTzQAMZcv
UiOG7iOqwUO8fR03q/pN48aooYG/cwxMUEyYQxwUhpDvqQ8D2mZSxtLUmlX42sBX
rU4HURZCFi3qbzOG/kxn1qmXf864X7Va+qiqorARswALM2CZrIchq0AHB0B4C/zV
mvUJh2mOD5+B7pwi0LFsQzYerILWhXoUo+y27M4oCvTRvrOyt2tz8tfYdrrOX6GC
FmOG8cqsp/2opGt28MvDrRMw29leY1egzQlc+ZUTu3o60lwNs7EgDkln1O3MNqeR
04IXm9UQPOm2VHLU0DBypan7/PsamcJr7IOVPd4oc0TF+j09kBJyUln34uyM2Em4
/CpowYxrRCTkyOc8ilW7krOpjs/u14ZNweSElRk6eey72JpXwyciYeq2RbHo32uB
vF8whSS+pc8bj49iU581WTQvoJw477wW5RRT2orXhIZDiKCc71zqyo9pqZrAH1rk
RRWXIzDwTqYGeD4Lf7K1WTPz00ap/vpvEyIWDd8+qRgimlKGyMLIm8vfPXUXGaIC
iiv77v3HZ2hdNYwhNcuisQ1UFAL6sHNPQC2Bf3GyyofZEsNAssS4mERVJdGdbsum
johm88tDTb5Au5IgZBe6aa/x1Kcq+MrfNFXxuTCV1CLsgGRidY8PT7qkPE4lI8jP
Le7hF8rkcwjzBH2sXnkRaO/bkkglzRxx11m7FfxklGvR+23T1ub6GMtMMRJlsMr4
G80tGBOcN/bXNaQfNW0g6ElhWReD8H+5Z9kW/GMP30jUMNufR/X4/ORL39AKtxjY
x73hmcWGF8D+J82K/ribHfji+gOtyonBanRmnjlwFuBW3qJs70kCge5x+g3/PVyG
/liyFuPnI8Hn6aR3qXDYQX6hlkmphhPWgUZAaFjYhceISV1I/MTrJ+LQ/KSu3s4g
SvtZvHOHPatJMMnFr9arX9PzAUUA/udhX/vYdA+LcE62RSDxQyPCjP7UiBu7ooZL
a3qplAMdgXSVfijPrCNJPSo1atDAiCdUnYNgiADuVf7/6apXbH0ouyGd12b5kiSA
AD+BLuk9AqAR7nMUGm/XheFFwe69n7IMcIb+jtQqoktJUU9nlIoXcgFGU+I2H5+G
emd5saZjmGA3dSlof7nk16Tax7w7osrgg028OgbcL4Y5/aUvi/zyFUCAkP67Klgp
WW3gRn8OZ0WhGFod+q5TVy1udPaCF1NhGE5htVk26zet4Cj4n+xxz9e0Jzh/rgv4
/igYoUQo9PnWSSD0MgKmLDJqB+PO5tqw9gZLpdX+JmyWlrfKt99w5Sceh2iEmK3j
vHQQq7qAQJ+aI3+SRBSjXhs5MkeNNvFUFuTmZwDqUTqf6G531QixJ9kIp9Pc677P
j01o73RZxe+fmCcWmrdY1etgQ0SKUV+v3nl/3qfHWzRBiT5kmuYbKiI2P0oXHKZy
EvZqy3/O2DVM114c5G2wnXq1cFdQJgjhHPQiHGwGZRap4evyxu9BHoWctFu7zlnE
vrW1jBPv5fg+mNkaaNDMOvsrnUGsxmewcLxg+rVLC7vf35Gqq7rakqKE1dX24yR9
g7pTWZwMjuoyitX7I88rP/K9wmTc/x3JhY4WwF3h3V9HW5LY1Z53csZkpeGsxHKV
oC/rteAn7PzoH7UpzBwkujI2odllwIQa0MZe/kTmuXY5eM57r23BYzS6puRZhx8C
zr/8nCLjOWJLSdpvV/DUpEY9ST+qWgwir9SCwm1sVwJdkPzivIUlpY6iHAeUHNGh
QftRCqzHCki3g0WG397uxWndX+ZldeMGs1C3pqM0LiphYqnG0bbSZkPC3OJiz3pa
7C4iaD+Kv6QvvHVlOpQBrQpszlkgcOKba5+Kvdauzy7IvhESaSUbMqTGysmNaa99
jm4fiMJlatUfl7BZKaNkYhW5WcRwr1pbk3DJpqxmY3iwzlZT4zG3y0XQqrAclDOW
tvtvjy6QLlep4oa7mbmMnk9mcuJeMGaPZT5Pey6qlizlwTaMfNjstacVQ1Omd5UM
tvFLzO5R261V+sSj5yWyyEZnXJhv+F5jshd1FtQ+ujabg2oH8TrYxRtux2b8hDTG
Y4HWENYLIhKw94oi448Q7t6BsQdwKNQBAellMAHt2rOXgPtzpD7CChHWPsJDh/6z
WQS8xGNtIVKBZsua733vDFlyuldfLTt8opLJDoOWtJCDgppwPM886G023TVXRsbo
ZgJkhBB4DjeinLehZd0F65VAZOWWVGMzikqaCS1wjjQV7g6iW6u3fvPyTPVXSEQZ
aolgU09EPMER1gItFxbqZg0eHK/NDlVMf6SLl0zyyu3qZHu2rZ0e5tEiO42geKCO
zfqNDK1iJ0sLPyBtsnvxlsaDm9X0nnSNOTVgS2wPZnOCghPMxMTq6gQHqSnVMXK6
zTZziPQToVnJconfgleJq8yQSyi+jd/BaKgCj5EpSjS0Wa1J/767K6zhKf3um/SH
OX9gP75f7SyrZD6nSfC0+ze3GfCIWMyl9lSpyyWXqNUxNRcRbmdUFLNRBi0tAC1Q
HBTViIBMDVFktlMdchJDWaStQPK5zURlWSJWL8oQwCcqB9c1T1ixObXMwS2lFYio
kM2vP7O9W+5CpPexe3fEMBS1aOp1q5Ftjpnbos2YheIDOt7XEDkd/MZl2Pc09Wjz
zgd/2uMnBq/VSu6bTKvIpLN5WobLCX6WXUV4Ym6iAg9WW4u4LWLzbaiohR2mdNOa
q8h4FWd4OKvo2mtqKZr1xUKV2xGAAXHCPzdkbASZ9ngJF9VTYEQVsqjKonhmy9Ro
hq88T84DjZi2xNWF6l/o8LfvjxrGaZbAgWUb2zJXCbJcpC74gehBs9T8zq/IcQf3
PahsaP57e/eUkXa7ppfj1N0s9w05rHkmlcQQ2j6/Zr+9pd3OokvXQIYMF5jjbEww
6MvvOHQCCDLffQUg7BpICcoFoqD0KBzMK3corZ+r0AR0+5uPp9xoGdWrlWl5vjrf
O07p0U5NjGQbnyG79E7OOLazeiF5OZwF2YP1FC0er28lP/EVWXc1xvKOCTqrnf/Z
8e+9DCE2NxlizubYJzsfr59BEvzFOo7K2pBc1ocgeH05MZXBnldWlcT6CdXSwZBD
BwVpk5P544tBTHBoLzxlkzTEO0o3ViK3ygIDH5H0lfg8JH3xIxMc8HE93BVK6Org
UDstOg6Vk1mXklxo9j4F9PlmIos3LN4J0yxCBfikixpbZwP/F4hup3EWQnkSdbSa
BO+AUT2VDw26CpyscOnm2c8uwLNtvC26PJnv0ZesXh9jIUnuWifceLeQ+hRermHv
GL1XWtj6bt3h5SXT1aSt5RoXwGMo1Rr3F3/fQJlkt3LTyvLEZfKbMzdQkpGxAEFB
B/KjeTIcoPnM8Uz7E8FtT7TPjw6gMYeaU2rxlfA8J44J2ILiv+qbd8uKo7afgU9w
jRTM7QydiRGaadSWd9cea/5PsSwimxowySryrfkmKlrheaql28H27f8ZkImwMZHD
K9T+bfFLjp9NAJkEyZGDgUlsRgKE9NVpudQYUYkk7/k6cZhuBYvTprTC1ED0ttwT
UuEFOVSMQHuyOTmLdeMUD/mGS5pYX4d3Gfo8d1ykgyIBsM788/hXz0nqu9UlATed
d33FhSNOPRo4kkSXOpnhtDt/p4WArjMhfpQu++o8fNCK0Jk2cdFsjcnBBbC/GZqM
1aKj6FxwFYp150bUGDAFPRdw+V1eYDskEKrpdwOhLWzO2p9KDftWlUbjb02LglQc
OvsJt8Omlb3+PPYRW22/wyUpb4n0qW2IzEHcs1+HPZFHP1vh4o0X9ko32/n5S7a+
9wSzpfrIgwu6t9kNPX0gtSxjFnXT7D1vmL6mrVnqNcJ06Tj0++OH81nCv+gkXHFv
rMRUiIAbhnyGQUI+lw2yCYuxoQmYOW4jcTrBnImacMjM43OgNp5YaVWqcvYqF2wO
/e7JRwOu9SnGnRXAuyhtnvBX1bmZJ1TmYffcC727CbWALE/NP8kzyWJ7MCPdy/cj
FlcDDPvmbeSBTQ2vqSrzEvY3z1LSlVQhUnwwAEzXIGrBFn1fU5+J0orjn18ludbG
U2iivKe68FlZeALhl7Qqn5oW9XDsskVCpqDKcViiLg2Laq3DZCGa8oxZV3qh1buD
ek1LZL0eZxQY4Y2MBoKx01HytNk8o/ijvYimyvBs0zddvokh5L60eFByPgPZlxI7
Rt0kKf9lfxJStxpV4gRkBqjaSrtbHjPohmtFMb16DEIux+DJ769GD5Z6D3LR74wN
XXmINPZ6yV6Dru1kGwxYrJHmqDAuUd9z4y+cFTNM04ZOJHjCgwL80FZHTVsvtFsB
FQ5Mb7yKrhLmRRzXhY9hTFGPCZQR3MhgUyNbVK1SuuLYWWJkvPLqg8Z2t54xpp6B
f4SeruGJN1xAdRl3mmV5T9sMbyv046EVoIq6AXydplg4SfuTx5bo36tJlAdKTg1n
KzCWEptwBymxYqAzlpuVV1nc8twC2uAlWCbjeYrLePBpMKRIVURYVD5C3IUO4Q0M
1I0Oxsx2UW+Fya8F8X2QFzN4A+yE1JBySBNKIT3B3UrtyGPlYxbIpckdDORncWkC
0s15/U30xlQIrI2Z4zJfkI6pzcCCkThMPj+vHsj9FXuwc7mrxwpLnKiGnB18KOat
rbC2Ep/0tAIuomROUVn259qKOOF8SUJsGtMrVTJGpRgwPrx6Fja/gYZ++Iw9lEC8
Qm1q3wt6rkHUmuyfDxxp+16nyYXU4pSLEh0GwBzzPRPO7MEch2RA/0nkLVWLvoR4
P6a20zCDI7ebCyeC7lYDjThVxeLtsb4MHXnMAbUNlpHinbpNtvZ0lrZrrGVu97h4
VXgeJ4H1WViXA4Skp6wjh+PN1FBDNQcCwlA9s9vpIuQHae9U3Zxiyi/oraAK+lOq
IRDpPi/iKAWHFZNgUmKmXppcsoR6GDdfMaSIzrI0uvREXfYrkazB417YYvBOfMl8
XQcCJLYtCv0OxKbtlRt0kfHTWE5PGI1KXvIuhRC/zEBui+Z9Drt/wNpVovZXAB1d
ifQUH3MGYOG85nHKfAodILiF4EV8H2WuD+WS3LzezkihiWvdFbSIst8NuXTvNQFm
AkIw1ViYPmkvQk9zW9zJzcxZyW8b9yXVSgza9FSUB1y3oEncNQJugjT5XOGdfMe/
4p5csfmkDZkY9+XYOuj27fG42MQQeyFA/FkVw3NzCvT0lW0X+RJESdvG0SCZz7ME
QZyCegIFvfirLOXCKfvDu120SSlr1E6vMlXXzwT46YGwAXf6bwTUerEPWTGEPBxD
QAUhAwVoABrbAW7ymhric4VgtMcN06RfqazYcy8W/gtueCAE9Fj+1UunNOfe9goc
M7IUH2TjTuhaaiEyQzO76o10QblWUQr/u15maXY8KQkDBanVYOyqXZYTEvWwWj6Q
T+A36yqmoj2DKjh7KZRvmsk2UXZ7BuSuLdDd4i17XnxjL1XsHrGbRaBCElZTpcLy
bj4ZFzC7QPSSDDYDjmEfuItxi19dNrDOaAk7DEQis3Q1dxKWnDi8GgYNvawjGp0U
p3JCF4clq8uhQOFhj+vsOq70DMoSxm2pkJW28RtvtdwbyotI9847ACV89/zxQh+5
qSfyrmbrkMa9WjwEclcGh3NbOpWRKP7s4pknui8vye1IOclABD7NdVf+YDvUXayt
8U2ejl8nYr2gOSWDXGj3SwOd5hxOvNFZLqnZeRbwt7kdAwTfaIE0kdcP7dH/38WB
Y94pKY5TYVgKhMS/OS8dNQsxUUTrbZkTeIuNL0TmU55PFWPm/4ZWJYPVbkzuoiTj
ZCKj5upecZZJwoqe7hatgYPcobRAeRrEmpcAwXKelQbSis6fPIsIHe8jaAca8xCO
5WQMkLY4uUuaKIyf5Ys0XDc5pNEt18zhIep0dT9cS5M/VnlrdcPa8KscNQ3pHQ2l
x1d6Q7BfK2Ig/TknSKhEc8eC6zVfvqDkdczwdm7uQYU3t8nQ7l96AxLejtE7nVR9
G7uX10ve9P+lX3VMUEXN6NGgzVqkJypLDjLlbo7hv67yVw35hVz0ByaTEemtqH04
0eigWZscqwV4eeaJp14VzX8UhMjJwOOtWHggAjD7jd4KsyL5Hn5VlpvB1bOGvhY3
IerQt1BR5R4yAlpTOiVi3kndK4nFzmaB0T5/vopSzV+k69n/+gQiOY+ZwWNqPvHm
e7zLfbQB0uMq7+V8eznqgR2MG8v4xJg/ruEEGkMl45mFZ1aK7fODl4wArgE4cmo/
iZMAL1KQvC/SOuPiUGoqKyUbTkSEHZbo5RPoQ6PQboTvlmuBFgj7a0jLN/jHhMxZ
OQIbwHux3YB69UtTM525k198Cj3m22rcBs6iAN7QYLWOJONZkVLNenemNQgsQ+Ml
PuV8z6BffUOAmJ7eEJs52QPv2vJHX2CtQ2TC3mZ856WWpswgO1QetD5IK081H4Iq
RrlxasT0dCiFVcEOuiDqyVPFesh0SrH6uK4iJnQ8U7ca2zey3XdyDXenDKxCf36u
dJ1uNmuVdVJREl/uGF0CQQmt8AFtci0JWkNv7VA0/dZoBwsYMIYybaOAbMdjrGEY
uejxr1HMdcLB558yBqboMBlBmmUV1+6Iid7YTW5IFprJXgFSCpdSPDg9no5XU/CG
0qojRdw1lUPfPL2zfjLeIV/BsDtdaqpHbfH+9hiiNTI2PEC3ZJ4Xcfcj9RWr9Pcg
dVNgH3X9Oz8LI4ZabP3XdwGF3e1AES1tSkKmKrwSbG12N2r+joTKBOZyxwmNhcQU
dBtzVuaJKyhdaIXmQYwR+Ug4przAQlRq0FQ8LWG86rVxA4UOlipEbjmV3sei4t0j
3LNYNkGeOjevrn1eHKefcXtNnagmf26SHD+IDTxuvbAKsvK6KE7siimFh2BzJGP1
AmjzKVmAsJWdhVJP6afkrOKFMsk0JuafMW7vkNz4QaUOY8DkqC1k8rhd8ADD6Xc2
RLz8Av4wzFW/BwYy2PkJJ6ZTWm27B91eeSxI81lCx3NAsXrvm32EJ3trDCI2L6M1
Pzo77afnLk20mdJ6BuMiTMONavpsu7gPT4/bs2Y1reiCTaSGH1f/go+KP6UM5mYN
ggZw28oW0Bq1EOOY/2TlrEwvS9eln2l8xE3+yZq0CKFlWRp0VUGf1SdVucCQBSF5
9lNxczOkCEIbPPbQAwTb+jGtlt9lCwO/gHWXkefqXGMA8czEapSDsUUxa3vJ0hv4
L14cA0F8Cy7h5lbtNTHhogRnLGMgKz2PSfQplVch2Ge2n632fFO7R+NSyddvwtbS
7NckjxrMbpivkomeM8mYShRjRXcnEyij7CtlZSeFYTSdOZl0h61+mpJnMun08oQC
NJo+JZhoChv+rHnajB7AoZy+J60ejTva77M0nnnw8I3A4MYD4upK4AXbKO58B5rD
dFSjxHhPsACV0eaIqy9In6aiA/CXBJzEmgGlG/oqXXfb/ZSs81OPnif8DzFK2Op5
lPwf3wVa1ZN+iY6KhIKDMZ3LqzwpvFwZv2qO/dIzDF4GcqMXB0TX5MrgT4ZNw6oe
KvHHRqw1oXVwF1a1HFG1MlFurns18z13FMTlgpGPICu2evjYJMOguoF5Y9+EzpLL
3r0wSFjs0DTIrbq65GzoR356FeCDhXc4hAcGSfuazUhMvClnLtEIFBxB6KWs2qHD
CYIaQ0fjgrTQw0dY9MSrRPB6q/rcUNfPgFIz4EpjxUmgubg54HvaOymR+osg7tqn
38ghsWXYOBrQz3tRdza5TS8IuIr/2trWxNe11rdaK8I0Ec5uN/yPFXU5qLQ0WQE9
2zO50JrS8U0v4od9JhzYxMuZOMkxp2/9X6YXPDGPRKjOaaBkGMpyjbYnpsO2+i7w
QQ03oaPyITSqSxm5V7Q9+GoRyAj0J7XYGLrb9lZOpl+uATefsmhPE+W7URbzE2qx
MZTjP2DWLxY7JQSOte8vA17DG4AhmplgfO0/ekvvyY/+SgYfrFhbFnqGIiCTf1ZX
oq/XX4ENDTKl1d8bu8Kso62kjnJ0mkd2CIAdWIcgKbNxxM1FpXKxWdt3aey0jSgM
ncCTFJ6BPH7ERwNTB0ozTthV5jUD0oYg+ev8OohsdJ4o+bdtfzrLH7EEuhyW+HV7
sLAt3tHOAqBCmQzVyx8C1++XQPhpYd9cFufp43cBvP2OqeNks5U5K/oAbLS8VxNw
33WcLEjHk2z0hoV84DasfwgoM1xk0MXHlka7wBhoLxufQW3NgBfFMmGFROwGBqHK
onal8dpVb24xLalr62Xu1AcVTeukXfiv5Ds8KbmW2+essscMx+N9avkovhKFF/IP
tpa9LgqurN4i44noqaYnHmDXWWlXcX+1Z0wCC8z3o3p+KzAR6+oYhk1Y3BThlds+
l3yzgBAIkjaUdGERvIWT102ymcNfcjerGSvrmbO3rEgoTfQZ87sq4E3zlBbonWFJ
5LKXFWuePS5JSrgDTXRD3tQDpeM+qDG9aHcFYTMrwo21GlkItaL2jd9VZC/jdX7g
OT/NK8PurC+XpgPX8YbEsgl4EdmzCl2XHdOli9kCnu/ZDrc3Wbkl059bxVtLp3Es
7NvzGFxFCmlebAL0iLIrSMY2LLMIYmnMiJqBUNROg6O2/tyHBu3n+uXdyFXkSwum
ZHyZWFeDpx1PLWeJ2a0iCOrGlgJPUZCGDsJnbi/FYRboGgBOtzdiMvniHTEUrA9C
loT/gWCyGva8dMaDuKIswIgFuka4DxuOwRb/kinwEgd1FnO0UuTHcPLzElBzEegn
8y1sjO+AUP+UWh4nAxZmoA==
//pragma protect end_data_block
//pragma protect digest_block
Hrc+yvDl1EukfevzMeHnT1l9SyQ=
//pragma protect end_digest_block
//pragma protect end_protected
