`ifdef FUNC
`define LAT_MAX 20
`define LAT_MIN 1
`endif
`ifdef PERF
`define LAT_MAX 20
`define LAT_MIN 1
`endif

module pseudo_DRAM_inst#(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=16, BURST_LEN=7) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface 
      // axi write address channel 
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [BURST_LEN-1:0]   awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------
   
      // axi write data channel 
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,
   
      // axi write response channel 
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master 
      input wire                  bready_s_inf,
      // -----------------------------
   
      // axi read address channel 
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [BURST_LEN-1:0]   arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------
   
      // axi read data channel 
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);
// Modify your "dat" in this directory path to initialized DRAM Value

parameter DRAM_p_r = "../00_TESTBED/DRAM/DRAM_inst.dat";
// Modify DRAM_R_LAT           for Initial Read Data Latency, 
//        DRAM_W_LAT           for Initial Write Data Latency
//        MAX_WAIT_READY_CYCLE for control the Upperlimit time to wait Response Ready Signal
//
//        reg [7:0] DRMA_r [0:4*64*1024-1] is the storage element in this simulation model

parameter DRAM_R_LAT = 1, DRAM_W_LAT =1, MAX_WAIT_READY_CYCLE=300;
reg	[7:0]	DRAM_r	[0:8191];   // addr from 00000000 to 000203FF

integer dram_r_lat;
parameter LAT_MAX = `LAT_MAX;
parameter LAT_MIN = `LAT_MIN;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
dw7C9jgN5kC9XYHhJu0eeNNlhHDHOoWBGOa4A3r05xOgyuFgdHg+lwC1a1I5BI0x
rtNY8R5TONM96+/cH87JSM3GIbuL/cTeUoebU5m1tFi3EjFbJxT22R8IEhfgAOWG
OhXLc9K4cb7vc5Ql85/GpXvCfJDRZkWDk1vjxkMXs04JonPIFD2q9A==
//pragma protect end_key_block
//pragma protect digest_block
Uz5C6o1UHsoLJLXMNK2xj9fMONQ=
//pragma protect end_digest_block
//pragma protect data_block
9NHAZGJCrqRg6HotlKTVsFKh4jBYLLhOaAGojpIV/C3Y9CdO/xaP7bAbmei1bqHn
sXKrtgrXndE5lEWzbZPmN1E/OgH9GfCQJNZ/xn/aAdql1NJHbnz99CtqRWGdYTjM
3WZEYAny8qiCcduN1j2YkAfBkrf6drtUGTYEct2PxhRV/e4+ErrZBBj2U+slHW3c
MTdxp43PiloL/fBekFe1ZWeS312+wrfEf6EyOHNprUr6OauXwxIo/jJpwyqUjjtB
NCQlYdsJa9h/oOjvVRP/QyXha6la+BPvVp7U3sl920Zib4gylFeAPgmV6mdoNjmb
m88z05Sb1Ykj6axt4Won7KwBz2YAFEyTzSIqxN260h6YLQIGMQUxe80DE9nQjRbo
d8DRPRJ8/v+yM7J9lvnbwa9foYj5IN+zaNQ5oOwMfUYDGNS9K/lBRwbrNSeiSm6Q
2YtOQHhw8hHLx5U166lxhozneM7Ls82E3wskixnu4DnocVfPiFMYyJQTYTELs6Rd
mXadJuyuOopi4inpotTIHO1/cwlzj96/rjLsnbMRCxCNIPvvC0g3tKquEUdL30uV
YSjrqCABOnOGVvO1VqNUjjQIDVnqpQ/0i9fTbauSTYIG/VqNmAxO4Q00VkTGJsWS
Emva7ylDdIyeiLmVxd38MSz3p4ptMOPZfUjuUupGYpmbU1Md3TNhJtkBDNxzGz6g
U+IP+Lpf+/QAkH+vmMMuJ8s9vmFrr7Y1KxwZ4yHZk6ExO2atgZYpbQSdH3q8qSna
KDlSp3+Zwo2YF8dwBruiK7SKteHZjU6Z8qhzZTKvTfVjOSTWB0tj8dY6ZEM2/Vp2
4QO69daKxEBy5qdU6+VkpZPaNSXyvyRo+XAj9y7AHQ+7+gaViHIT5cz9fyc6ewNb
WpX51qtbHD0i8ELyOFKNiya5u4m3GEvMR/jKgtTRr34sWJNYVfpqawVUXufBTWC0
dRWaUOo74DN3NnmJ2LnnC+2GiaSXnQSGvUhGCQ+of2L3YaW1jYeCB0PkDLmnznxg
aMS4M1UeImPt+3p5+tPzqFe3IkrNNWdQtaKU0DXyId+ESFgqBM1b12w33/PIJipK
+zlrkVESmcDKWI2JUDQU60gatxLo/HFC8n4CVChZmnedOqMsCE1XFKyc5rFSgkib
VQSG5ndjtxZ1S0dZBY+tlPizf+DAyqoD5RedI2dK2bmFlO33oZk8MGjwzB0cRRnH
HkpRQO5+wckiYiYta31xnCgWpPZHcE+A0AXx2BSNVE9Kk4Vw88IHoj0Ro9jtfMoK
fbuIU9kcF95lLGyGdLv37ooggxb5gLHVAPsba1ymVlugYXZgl4vVxhfmToDOzJNn
3gDpDCFqkhePOGy9CLl7HSepRUizLGQjPb3OtZ/kYYbw7zMK7g8wR1okQPaFO/ME
hrGZ9zh57VxZl4Wbps4BHM+cbKd2N6aELV7Z8fvWgRPbbS18r6WA01LAGpnlMGCx
SQRLz0CfSvaALCjXs7aYPkStjBDdK57oFfObDBhTKiBqALcQSn9aK7dnC1SuMJz2
z/L2NyGaHTz0WGcAyQJVW9rd+sUbnD9sqGl1+8Xvtbht2QKdlIJ8FcGjDAxT1Zh9
1nlxef4MlXrj9TgNy/cvyR/85Z5+b7Q9ELTXl5Nny3dY1MSftOEZ8C9rF1+CtQVU
Y+9IfgZNB5axNYrmKBXTJethtnGhR/ZtsWP/0w61WwyDNCoM2Afk90H5MndcZsEg
Wm8gZ3yy7lQbws24i+Cr4j/1sAXo+gtsSJd16dRuP6tyPUN28tb1o0S6Midfr7f2
gzWfBM1v8TRuIq30M/IH1yQK4VmaArRyi7LtjSlV7lfDPkBjCLJOV9Q0FXZk+oXJ
gROcvNHiQ6Y9JuNtn8indvrFHpVMErKaEfRhtvb8tGgAkQLjPSoBuQv4xGXh7nB0
1IaMWs7tjh+SBwDxZpCxrepI2hGb9okH0Mkq1u2hIuFX+Y32M1HFHAoy3/FAKOt4
65cMe3RInEcu/5HAr1ORT6iqWe5r5AeUHon4vpUqcdRm0buW1lzj5PRZcQmWAZPh
/x1c+XuBX8N7s9XoCtHVQRFjwlBlCSogpcfpTRwUuySyLcOj1fs5loZS5bP7qAfb
v6u9mnRfdi4m4NVfLeZueeHHMcDi11tlh/0Coczqz2EpheprJe9xKX9m6oVPv470
PY/Ajwdwt8ytVij2pfxPHw3nTfMtyY0VResWrNppYRvmDPtSdw31lm2WyEgya6jb
MlcKGXZV6x2YoHUlVH/bVGOGVTAMl1TSbrbH/mD/kqROYPmRYTzHKEFixcl5SUhT
CGxMvTgnilbSepFizvxwlf362U3sW4pgL7vwyqIjhyexrhziMVcS9CPOgmXdyvm6
adAhLDqTJIA3RCc2bhctue0mF7MMznZXRq1kVMKYfNFIRtgH0n3K4JFFwJ9B+UVL
JyhdDKEB3lecx9/kyLUGE8LBb1OtsZrbPfR5UUosztzK80a3U9quNMLd+2hbwGFP
K0IwwZkkdKt1WLrtJMppiG6oTJftZOtKP1F6qov+rob4EdY/5pbR73K/+yYsdIvr
hdMHL/CKQaqMzH3HGhhpPpGLTc7FQAV2gN2mX2nOwD3UL9fEqYhN+veAqBmw7q4J
Iv5LUUwqYXwAy0QsOstUFQk98I+H4a/IlRbd1FQKxiu32GYc1mmilg14cKQa/yiv
SPoI70GLbpNtWjwJVwy+2eK7NgCVzQDC4Pfh8gV2tQN1hhdQwClFmII/+KNnsXEQ
AlNXXUj3oejMLC6bhdAJxKxPpwKlx62toDut8QWjF1aC+PR6xaxCgqvKk7jFByKA
cjHV0XiTBWBQtTSUnxa7wi41bz6ETaWy+516L0p0J5KTUWKlxir1jTH1Ug1Gya0n
tuBTJ5xbjBcvt2JAWZ0RpTPXGHGRI2C89OFPe/kDHIjHRBCJ2/zCnhCgK5gyWJhQ
9SxuN9ZTnYY2T6+tjYhxUuJmkgZDumTTmu9fsV4zBCeYeWWFGv4BWsAFS2GMzMoJ
LIfKdKWUwl/PWZ7q+e0HtpHUrLWABvx3G7pbM8dtqSbSG3Hjf84UFT6AvV4sZgc6
w/c1FAb9k9vNW6tuUdtdxkvIsROYriLYvRWv8A9f7ZQ15H+NHtSySHKlHaHf6kb3
TOUIceSDeog62/coamn/ICUnCjh2LFOj4JpurMcbhFjuPIq+6LFDrb/WQtHkdsrH
/NAvkdj0+PvuX7gx3Ive5dSJwPJlss38hHb4sTx9wOg5Q6S3wuGpeapCBPesl2fX
Ose15L1niGhjX/4gme7XGMgRMZbmxKJvT2B3VaZmd7Ud/rveIUUyNomDUGkTX4Ai
Wdr1bRvVhYKI30wuE6sHnpm587wkNXPsWVY6XB2RMe30WwBZ2CruUQh0gUHRtqdR
BdurcgDTGgjq4UdaCTFI1mZOfeIgPHDK8wfL4U6cewL6PCIsLijouTB+o2pqeILY
jD96wdMNtLtc7t6GaloLu1QwYcZOKfuF4NiXIQNKf2A93HBiWFQCZyHMulqdL1Pb
iHLqQE6qBhIILsj5+SxHIewj25FGl8WyspVIYwSpxzJUQ/A4ljuzmEb6B151fvDj
wm0vFp3PuIEK0Gr1nBVPbvVp4JDsQnhhUBUghokqOiSlbiYif5tMLESTzSwE6TCB
Ket2BVE23qaAYVQKB3pH8A9p+qRTgYf/6ZyVAISOOWoLv6i2T8+40Zs2ONIB9QSX
t8dwdyOva+JUD1U17akLRCHwRatIQrhT3SyIsETL66brBbP8KE8UKTg+zdXgrS2c
1GT8n4cROKPaOIVkFGJcPNj/MXJg/FcAwa67OVqRw8cd17fB7D3kcsINI+2Ok/9Y
eTgvDhqUuBOWWA8itrrvktawVcJkpoXwo0NMd0tmFqGhisQ3zkRUBUNy+4zf/cHS
/p8aooWfRDxxcUsvx/LjTBXYSccDAc9uXrtFgsqfr7H/pMiGwYG+XyrCEliHcFQt
Ua5I1FRDiq4jbmF7MsLS51E5cCBTrgHZIc/2FFnm9IAlTGa10xxlepcuLIlvxYaE
qjqnhkDiubrvZ0hhGjykDXmTyfPFo0IqwPZKqfdPT1HDFc79SuCu2iETgJjClFbL
SmtyXa71thA9FYLeFyCfO4QBxUN1OYfabIeGSbaAi7Vv/2QfA8Mrr8mFqmBivvSK
0v3kiuUFiXyQ0yd8VC/i5GYk/od0UE652H6QMod0SZIl9uaxvHTM0WZMiz7oe3sw
7VT1AOGA2dfJCagmIA6VJE+gguuYxGmyOKlgE9xvuPrxj6PLPIYhgHqzYfLrFZ0E
rSBOkmD4M6ygReZNTaUGF0X4SiJ10WH5PkXfQLJCw75ungUxevqv63wXQ+KKFfRY
b78Om5UWVIF0fqVIX7COEK25T8NFiBHdxY0Ea0JiVfXT7at3Nkpcp7+6NQMDvD4F
HRchgygnzi38UlbN9pYdTOAW/v2b00x8iaWzJYCKzW9CqWyxADfq0/n4/tR/hIVU
ItJcDzn5P9Mkx6LPMOJsw+I618MVzByv+jpcHK3vuhWssIOxNinROZO7cBwizptT
LdxRKJKUqLOmo1lkouBlkQIKZLLC+ChYG+ae13ti2SFWkDJLKEzYvYUFYz7pFNyg
PTrpkNSUx+Tjo/Q/zgdGt2+UjIrmmAUg502yn8CEaxOz4ICngE2Mej9jWoaaN9ay
+MjXl9/ExDWO2zix2sWtrvdEDZUoLEQI/cWc0wY4GUyR00TPF0Xj6YWLDa3ehnP2
TshUOMjwZ/uBExyGRndM7r90i2IG6BwxlP+k9PBlnOBV8Uaz3kdvFUPD53da4o/1
y+v5y6LxKIiMYgMGlQBk/B7bR8YFVttuPnfTh2TsHE8tKw9xduNURr1rN/TcJJ2g
vxdd3+zDHcWljEMDQNpHAxD1SPN9mjYO4hvJ/wtF07Lt7shQZFsZ6ow3iQqTXiPH
D7FKCZ2U29QZY87T0RlAreHgwE1yZdJaJQ23qVEk1im+i7E5UuW9opV9KHdji2OR
wPEgjlHomycJye6vLBJI/P+lJE1splo4xOopCGWtMRXGIyxZ+dS6kytY/FHdjens
JT9GztU3rcE9RBHmzBAczauQ3/tuDGCk+kMTmnIFE3jQkK5MEFdHfUQMvqP4YtDb
SYUOY6ezrBy1QlZwVkkujpVxRC8FbBpIJBnG/JcZAoAJqLcUZHxKU+hLl/NEf5rR
x+q1eB0EbC8fwXrCvwjj1dbiNWJFcQAyijw2gx8cU6D6fymLjZ+xF30tYEq+LPci
HlHB+x2IRhiXr3FOSYFSyzDQPIZNHWTJmVd05Z4fUrhFdhXZ6jtaLp1k6ajaFUj8
nzqH9sbvIn7uJCP2NKKjw0NPFf5yJND3p7cVy0UfXqOT1+fM/DK3XQQC7bZYbNGl
Zpo+ipMEP3oADt5Iz1emzt4BhIXTJjl1UsDd8sazItopyioflV0Ang8VmwexJwHa
bvBc3s2XdH+PDGqZtTt4zpDnNcdR3TygfPP1RKQHRpRIwIw8+8ixscyQ8PE0TLH7
oYxIY6RJwKqYaW0f76wLjdSDhaWM9Kfz6xKMl1Hqe95pKUu9+ENFNbHypycLgMj5
uvn8vh8ByBJuYSe8Hcy/UYu8xTPgb8PAqJ8mdL7MBkwvdNCNR/yc+EGB1/SF8WBh
0Jx1K910Uow25vrqJhFa6pgupqQBHtoHtiKKjF7yWIyl6n8hxidA3bQzoz7X2c9t
HiVfUFOuhtNoRoQWlSa6Oo1Uyqc1P2tSzUt3HwGI7UmNue9h2oOp9NUWaf03BWgt
KQtG9UFLaLLExBTuhLpUDRDFhzHpmZDQnBTNJsbsf5LExrMPkJ3u1GndBC/hKeRn
GTxKupr1gUAttXIpYwPcpIrl3KIBLoQHagsYWvf/7Znep6JhL+jZFNb1JpuLnqLS
T4piVneZrxCqW+Eb+SNHe0wVk9070to2evOaDVocZJeWo0xpJjsgwnqcEchw2VNL
uTpeYnzoPL4CPhtnRsFyUcyVAiY3qN6uUk7gcnmrCy5E53XX+e+yb2r2k6+QJC6t
o3v0uL+iAY3wJJcyAuV5fyKNd276paEIgymZuGcL1qMYrff1I1JyVT6fF+9kZsFi
VdR3dbrNHWnhpiSEMAAlHRCYqIt7AVxlZDmY8SKUvp2/Px4yq503MHY3VasLCltd
DwnVjBTDrYZLZcFHlugLcAfLEm4LVwhx5msIOAQTTFZmHyh38iey9ZPCo6jwNyyf
LRd4Qc98o+uGJnOIrco0J+oC4sGoRW033x0dJmXtSty0UF2r7+iuUViYULjSzH7R
Ew9Wy7eimKr6qZblJ4kiBcUVM8pyY1tjLftIBSgdoSkTewIZW3quh3xRgo7DYkv4
idAiSRrjlMavfXquTnOOjjpPqfyGTtx3FznL2bWWE7Ji9F4T/D4p5BgU+LcqoY2y
QdguucPNva4FMsojXwzLDCnZGZrzBNVV2LlpaJtzuJckZSr4lNzn97Hc4KdpJEml
7zponl8hBWgp1dcij0ZUIGyfujg9oQ1xvxVHpXs4z9zfgeZiHINV9ax+mt3nyrn+
da+USn2VOiSPpgtDpf6F6M6ZRsRIcH8aB9QvdjDDmD87F/e+CtTg0NaJeJnanb6k
2bxJ0be7MtTbhS0GDrhg/f9aJLu7gGaEhXQXzzv7ASTahHWI5+4LnKl5JHTxX55K
YFvTzyb+mOMucyXQ7aZhqjqediizb2OZBzBcdc3t3ti0kYC+16tKbXIRMMpY19WF
1b9ZlT6uLkmetkIg2az0x4HeNpTl3bwZJnHNGv3BIj/A+zdiB2qDv5FGniBTt7YE
WNLKprAaWwQiBjVEbir4snu3w0om/ySLaCQ3Uy3HiGJlpYg9sCKuPVpnzcWabTvJ
w5XobvcBOeRuAEhI3zhkr1Tx9cGmDCwsKKCmPP/ut3T4K9GsdmJsKiWVOZdkWqp9
6dHsGuPAPuyROlV2x/ZGlHFSAAJ4wwACpI0SGKzCHJsOJo5aoYCUWlUutCn8kGBI
thQPBtbHNa3PlAzpSsvGw1GclL4h42ykJgIjXW7V9Fv7/zSb1XMbDTyMmSkF6meK
3RA89f3yMY+V6trGOXIRExowY4D0U4hQf0Sy4crtw9wXmHILzs/IZhE24DUpqWp1
qYENrJF2qNRa4mmdiBfzf7V1PdAKUtwju6RJH8/S25iu8gM6d+HuRpLkkhK3KYPi
LuYL6wXvDtPfHikl07P8UhHqZG37onsGE9JGlmisxqwGeB/WEM5iSwsHg1NiuULg
CYE5uNRntQEv1q1XcHXW9y51RnwARAiNUgvTM082wX1wA+EpWSHq+wkcGmmNWRqq
HKqAsaHab7qvMPkrYGhfQVIS1eAdVwFeDsV25uo12tEhos9Gp8Lv5tUdflUCS/rP
X4ybsKMrEp42JsMwKmPF5GP2BraaY5Uo5N0YSKwWuaF+zXYm5nlyM5j79lcq1OM0
7DK1JVF1U8V+BqQa6KQeOhVHRhs6lGRbNDAWin4FDPSTAw2pKX0j0sZ9nmHaqvFm
nEZA+275PSDTV/d8tB6rIfQmneDOExZtHh+Ae2Jy3SFSrM47rp70PbA9xtoDgXx1
fjOTYz5pWQmeOdfklhUAapLmbicqRpmEgEv9cIbFVREFlilDVwkzJlzIcFjBIfip
LqOSeaFEqUvR9ZRaNjgujF6IZEG3/0vgJ8XAG2E1qVeOtYl8WsPwtp9nvngz/iHk
zdYHZdpINDE5KMnbMKYUvDKy59ZY2OTFr3BB0DsXDqmkU1Qn3FXTbRPX5BG4P09Q
CwXnoC1SVtlz5tCKSPwYU2cNTBs21Ze6Fu3A1mDX9lcX29BM+W+I+pvtsHnAk2Vs
cAo2FB8HBfnivZX4V5uiBBfoTrnKnrjThPzIosQuikKvPo1dQR0ChoA7ocrvhjaD
RClB15RwFuJy1eFLIuH8heEpKwR4z8sBRRMzVknNkJluET/BoYAIb4xm/z+x2NOR
L72bT3he0jYq2g9wToxIDkUdmXVyTe759FD+/YnpLO5cMJh+1yVc0FdIqu/tsj74
MmpPJ2do2z618D9quhcboReJjx+F8pNmvaCe0Hl1qk9virb1+h1D5nQESfT7UhjC
4gmiDo0fjfBw5VlsZzaDY5sxDMwolmyh7oeFQQPdnRNwD3mWq4ARUQBPivXPvnU1
cfcfZyqdsZneV11kz+F6O2s3VvVdjWjpdFks93wqg6YAkp01Q4e2oxxchDkyonYT
SdO5G62b91oCV0Z/eVOCzTf9+tlYeICWCAjigyglsx0g0oMcRgQ8W9TYezqVADEw
aoB5r44C1sJndjRD0NNfu57Zjon68yDWY4IkTlY40mREcU0bb0u357dWqdCCbYg/
WH5ln4O95tmRBZ1Ub0Dw5khTQ0sOQRWE3o4TniVyG5CHlbmTL12iiAxVWNKGjAgY
qlUMKWQjnzSoiZPeXGqtMpDMdJyYh7UKoAZOm22vmezYp1wyUix0zKytKkgjCHwR
K/hH5MVWw6iLmO1HH+7Z0iCBT97egQGZ8ac6CEH532vfwXaxck/MxLAdVEfBR8gw
LwXgxNf6ZJsCfbov/fvhZHfnpzfD/nEYbCIIO5GcCZdxSaab4/d7dg7gwnXwpL2M
jdXONJrYE0eSbHko5F3uEEUxGqB860yZ8zQMxkR/9aGvJIs9Gu6wFCI0rU3vhKCm
pl0VbTrYr1rkUyzxiwWZQkzFD55t/bDBVWxA1WYxCWHs8kerFIVzW1peWuJzwuOQ
FJ/B55Qz/V5gWt2eR3h+sTrUDdhbJlxyoshbDmnUFI+sHohRCzkjy4Ojd1fmiOzy
xybGo85bVQd6VhV+v1q6ctqphYFCDDpshk+IAFD+T+6mLqO5XHehNxV+fi84p+Al
Ez8e8dX1XPO529dzlbjJCoSSWKJODxyHzOFBpE8MCu3V4RIvAHsCQ6L2C5FSMbgM
HZABhNvBtY+VLYv+IaYMEKjtdj+WJbX+RKRqaHwBgfXysBFuPUr+tuz5EweffCCr
bVx1FQUFe8UWJblQ0QMCFpFj84V3XK+orGWaFE6Ngw/dsMFF7DmHrk43W5Amd6nL
MbtNGE6Iy4dO/QKGXakXuQmgQQXHW1K11dU+VFiUHcCPjmISAigc50IUHKofxU9v
rOo232Mm2cgMNpkH+TgySIl0HZ/TGA8qhbddRmS1zDWC0P1uM8wp2CaYf22hW6N3
dPU8eal1TzWV6rSUp7TqypAs0c7hBlCee2awoSACYcP1mzieGb4norZNmEFf/7gw
PXo+S7iiHnNbnvfBuic3tT3lO/rSlkccjO7J3XR6Qo09MREUIKLZKQDHCXlem8lr
BVY3f6PmnxGJYrBIrLSxF241cNyAGJsRsjwVRc00oKJV9VPgr/D5all0HTme4d4P
9/il/nRCjHUCQMrSHmNYPKHWVGSQnXc1vayHDRsw97lio9kADPVT/UKGAsg76/mJ
EUCZEj92SElTMgUwL2Q5+/2FNg1DsytWDbiSEmqVwfsmUSgtRp/qmOuvO0HcMki2
q82OByCPOryOmWEqDSb+dJM+b1TfdzrKqmvsVyZA6rDXwF7S+oVJcjeIvTzb6r1D
7wfOGAjefxGkZDinLPBsP88jgMJTWq5ANddmEmuS7dIP0W26mLlJEw3YvxoU0rr8
ehO/wrdTHoi9LTvm1q2+rRLZD4iv3Y0rWIGrIFV9IaiD9JE+haHDtz/G7UFKXe5I
7K7XJzenSp/xs4JAmZHEekTWZTXYn9tQ0LCsKW86k/C1Otll7IwnyfAhG11AHraF
fwcVvh4ceESk1wdjk2EDcQtYjlS0WbTkpqH9yDo5rHWbs2P9ABUh2QDL4yspbRmB
owXEmDeNEH57V8zffCYPMjpbZR86IfOayvMIMePCR0ZO7BK93+XFcZzDfbs3MWPV
6QHGYzdlU3VO6k8roTHKrxrGyDyTdCoFyteAK1n/qQuD6MZ3Qfd8FX8fsrHmPQvc
1ESRKexnwxjmHTQUbbT8haAe4F/sm1kqW74m8Qd23ZTU1ScwxUGAhzkeTB+f3w58
UAoY9bjLqvMBUKus7XvPqFF4GYqUSSseqHUy+L/7TQXAPZ+6c5JTbH2aFwpy0Sp6
8a3fIHpNB0JvDi82k0hRybxNoV9Av5shaGcy9mtZE8qmbg4iiDG9ucOBiHBYLsb6
Z1m/XJaLedOB3PZ5jCY43IMTSzh7hYrZMee3ac/gaq74Hxu4gvyA2Pact9oVrMlE
hFZNjdMpo7kau0P7Als/CVWxKFBqmqanNn68e0tgOVcofMy8j3vcnatlraaEP0+J
I2+O3E2H705tTGH+zxLYEkel7wVJrIakgGDIn6ZaE2b4d19yjAbuXkL5IYS0f2cs
xucXxbDM6BxQOo1f2jJGUoCkVMO3ncsVJ03T9GyCqP2568plyL4ZbH4hMzMz4pld
aw2xwjZaGLhy39zna5Hzz4gGIoDg91Imb+tmTpFGBs/xYl3ZgpggM+CzS8BQp5+n
7dUGoLowhdvzgVc72A8eYH5/xVym/BOcQwLZEOOWH8qKzOceTkgXohhQFx4o6cA1
WEeCeXqvhSIWaefRIE63sZ3iIiLijs4gSdIkJz/pXWTF8DuNVC4JoSo86GqDX5uS
6gptrwyUkpLzPI2XgdYL23lDQFCTulu7uI5pysR3gCNKX/+y4yn3arUqvWrnkXoR
DE9bOcrzqYIt4aoe06srpuycgOHM8rZ2koLqfaJUcTz+qDhJkwFt2vmpjC91Ntbh
0w32wedGewq0eMg73ojPL2Hm/iiQfyfndQcEBQXl4/fgXBadmnrbVo6LMVrTzd48
dn63b4fiXZ9Alsp7duN6tMZo2rDwW16ACQGyeWFMv45cBD3rRhI/1LY3KglC5Lsv
H/EDBFxBd81VO6JiDRbXRMjHu6iamVMRnlQNZXoZAdahSu9ejo0XkRfJG9HVVxNE
bx9+lB+//QAVLId6qLGRjFDpQAYf38ob7uC0TDMgzKwjUnLlS/zY2oQOVq8yL+/H
k9EIwLLOECdcXpxP5OkpRKdRuuenMTsBxhqziL9Pxmlqbiq6h87mKqkbt7hAvktn
pZTgnzvx7kSnkT7MhY8FR8ftMDNxX7+vTBjqaLo7lJPH7jFuxX9q1tvOCXiI8B2q
rkXQz8JTwOBms0Mfrn+vE8ZMbDRdC+iezr/AGgePdu5uatcoFYF9oV57yvIWQqEz
X7un9xqEetTefmMQxmxq7uPKVZszWHHaTFlo3I+0cFan710D+groSOwq1GEM7+b5
YmDAJlU9O+Oq9iLcA5rk0dI6+e49oAjk+Gs6Dy6F1gN4EaOJm6Pf0QADX5lH5gZ9
xGqvr7zuO2jGwTKBMLN2oAox2cg13eK+yHj7pGcqmYftGm825YwldRnBxnGCpeZ4
r1wzBwZ2wCoF1QG33ZYAHgzYC3jGkYUVdQEu6Gw5gHSuFvFJGtClc31GXztCHgwh
mBmkj67SrsnKBWwRswXpdQfXCfnn6cjbQfUN82Sju6JSJrz1Om6ZtZjTWpGwER5C
eLAdgGHryF5Hd9pKfoDzCu7vyrmlyctIrl9ldHrfrO5JPC81CM3+i/+sfwV904I9
x8XtU0XkDM9RWQQwzfc/NVbnNU3MmAQs+yKG+LE0fFmHvwNoohIlCgN09E+QX8XY
eNESutA7Y1Nb/20OAanOF+SthBHOBbDlJ+gf4fSyi/Hv6LfpiKt1P5lETDikqPDD
Sxtx9MAHFYIP8cNjWk6WSB+5ofRTWRtGy0/y7k01fn7HiBq4ZbphDq6xHn//KVn1
dHtVtlfh2eJ2nO5PPjUYUtpqT/qsLxcB6xYOTEw8V3qYkZ3DUk5Xgw399QAiI7yQ
Jw6qiFVpUBxAQZAcK8KYMRq2xvaaHcIAHpvaNQypPT9RJ4IsOU7iF3arEG/KTNe9
pzv/MU9o1pBnzF1LlSnYqER/UsLzHii6j5hYIPoZV7csD0AzE7qorq+Yq2lPweC2
MDeSPitLFgpWNiUEwIhFdZkSNky41cWfli8yseshYO6xaTOfeeINNcQRdE3dsadJ
yHAtTqbsC3EjiJvrZ6ljhvv5gheBgNJUMZeUYAvf/DIgLlvqiG2rXjIXAQ7TiJSq
HpbCjESRy81/YnBf8MLvk6X2VnFzWjJQy2/5Ute/Kkt/WcvM98nhgiszGHPnEu9/
5kzfELS6h0vM9d78lcJI7Nz0Ut4ggMmV2+aIDTptdMCpeXM5TVtggd4uuBKhserr
M2Bxel42cbapi+MWbQpF6vhlFRSpuOw4L7FIu9mPKOxXZW0BtN5pp8E2kZGMqs1A
HmUevt3KSk8v3tp4opGVwHYjf1K6brsf6RWuVqzkOh1xOpNzODucILk+ZKDXlcJ0
/ZIABwKDHAttf/bG0R8PpGQKL7arS+uuZGGRGtVqWL7uRW9rpmdAaDusC+dmcoMc
j2TOFsWLcbA8e6+SiaMpfDnZPoU7Lr8ueDCE9s/OJ551cacNwqJWBvX5HYjvzaqd
EOeizV095/pEvpKUhetl7B1IWor/3KVBO+XF2IvRyFIeEjNeUpA+pw18M10zMX2p
T2NpFqvzB3CidG2tfCHGt43hZuQ7GOpxCxFGpLzN1oI768ZCVi3PDat+NYhi82FA
M/iQKz+7kvaMPLy6uIVD2HH+hJeTJrBUTf+meuMa9LmvL1h+1YVqCHNIHJn/27k1
uimSOxi7vK3TS8LED3UpSqy5q7nOaAmRkyTIPy80+opWuo+yRMhOCnv6paf8dTuy
fKB0Lm69PM6f8W9HrolbUuZTIFgP1y1fWPC5MvljU050bMPhPVL4UzIcQ3e2sNH/
Lr01S/9Th7Lp0hj7bi7G6dYf4IgWHt6f1c51Q+28j9Te9QKP+LfMQvvRfdbZnrZE
uETHrKJZwiQ1/DOw/3yQDle6QD7CHGu5hEu4Ffwryh79txEwP/wMtv/bDeQudGqN
Fm1T1X/xVSSNwa0muzOhMiYv1M0McdPfJs1O4hfVXeQ7IiOTa+TaBrI8DzDejzpB
THcFd7ZVd/87qm78i7C+seTifZlFT7la5/SOvGeSXP+HYtkRxEF/J+YX+87Uq5pq
7wdiz7wNB4ZjFyBVvl1dxroSFNodEsOUuGtC0FK2V4IXS/FH9CDLvXhJ6972di6Q
Ke+jCmPzgk8L7rni5tBL1HVZMTFvYJ2Zh9fIA/N3vJaIravRvONuUnB4dUOK7S94
0NfQVqM5ay5XuboKcl/tsmC0E2wEnIYW6t3e+3900lsV0WnUAFh815QXGHub2iVI
p+dM9K9XnsLPgJZHZ7wf9teqMmavNCZEd0tLaHeHRhLB5P9pq3B38Ve/CQVFtBYo
HrDTlGe6NHIPSireHipvXwvHYn9Uh/SOsUVYvh3KvUgckOIhv8yg+aT4x0CpjoZ0
nz3/7FOoN4rBtAyeGzIK8xRXyqFrh0M36n/pyc7rqlKWx+O8aufM+cTTorFcNkc2
pswBP9PIovxiY+Ytkbtu7fkfDZ+3COQ156iT6hDNYIDxd1JlcrR3cVYBrG4mHBxJ
N3TGRy8E0WV5kmv4q1iNHpTK6xFgY8+xE5wkZNf6p3TqgznQ0u5+pXzRhMYTs6+N
x725JVwGAxI21giakY11D4Ol6Ya+5wwycQ6Y6IHjW8bJVL8ybbfjwr379uXAeyFL
ROAJRzJjbzJpqQiCFsVkxZMgSMX7iFgn3V0JnKoiXj3fAsLBR1rRcCnVU9N5uTx3
16/P1Hs56fXDBkIDtMWB8mC3eEAimYx5SPrA1HUxksM9uopvYFlJnxzw+COZPY8H
TGZacBZwofzTrVeadki53oSB6airQjLkrUGRnQe2lMAkABaqKmag7SvTPwqQCYmc
w7ypw19j/665EBxgE6gobq504aTyMvrKK0WneCJX4NB31mobVy6ME2pCGgqmdLDK
DruXfShUGbuaAN/yqSAEvmxpc1/XupROb4uAfAbdFWheOi5PYH0wScKxMol+sIaP
VbtMR5t6S/ecI7YgF8fFkzdLLmch5ylCRurJeQHDsG8OtcrXrGE/vXt+PGwXrDRF
EeC/S+ybhPu94Y5ezbf9BDqyuW3F1AqjKd5apXf4ADeZKp5/Zzev59rxu6lDGCop
OlpfB8s4BICo/aI67jfaSW+XNOdEc5uHhLMvL6ih8rnfWrrLdudAiLSN+RlYjmc2
QhQP+rF4Xlh2IX1oDnWv7lpajnEWbxAWaDgkOf4V4ZLjSAYXjcKQV9kgwhNkqcGu
iW7bzT8kPalLidmrhBfEcDNdGztQVY9q4qgCXoUZprQddIhotao/XHcfrJr1p8TZ
GkSm1JWBl1AvbXb4wXWe1U04exvLXeq967SIPntebw7MY3kBDEFAKgwU/xIhivu7
+EjQQVzGCcrnnMvtDxK6NPe5IAxaN6hMWkhU2yWg8VLBAu7oOzSSroL9GyNaYBc1
KC4VrISSZQ0Jyzx/++2mhQl/hSANz/f7t2eLxkAQA9mCoe1MOhlG/WpZUWUdvaH/
gkDOHwsA17zyCAG0rdNeH7BunGvrCwoYcZ74KmzTi9KWkWzYmhJ3tff+kFBkEop7
eJ+uHGGp9fgvctrnoDfBaNkOlUpoD0AJE70d03WY2TXbXVzP1J2BjdIAkyaQTD2K
LBGFIArFCXC7VuVAaKbNDcm9m3KrQuPVq+bCEVQAecxhjdA/VjCLIVB6AK82tbLq
5IxJ4em+vxzIip8Zq1c79SU1JRD6wVwCpVOc43QODCfrtlA5Kn5B5dNtm/4H0mnz
PqcrSSNXHz1kWfYtPBgAXOk+lgVhiL8murVTGVrtZPZF8JnkylvA4VZzcboGfRAd
ZUKb/Wr0br7Avs+OWluCBZty9PKcRbW3VyUgqs9vmAmEcVZTNGGF5Fh5csYZw2T2
dwQUQBFfZiUUnCBr72Yx+HDNOnwSVeqfjAB39aEsyScpVQm4/B6Yl/HCH0wQ4APU
nGlXy52VbTUsTpY48Bt8cgYfgdslfnHZtrBQmpA1Bq/vLBb7XfKxjMfpGr637dGr
wsfptkq0BzY2RfBHt6YatOvKRp0uRrmGk1+uB6eSwUTB9j0gQmBc9S3tlryUsmq7
51FlrzVegY0h2jxk45qGRSiOnvqUpZd0ypZkafyCx8mpn2qUQaOavIDCML/YZttM
i1HN5fppMfvMsuZOcioKyHbgy1ce8RNzJA4PjoAEmzpCHAGgBBOZNRIdFR9t0k4B
/r48Ip9qPke+2QwlScXIGkoawzyXiv1pTJAbvY+qZgLe2ZxZKFF3TzuiD/rbwB77
9RzW5qtBYa7y5J2wDlhvIXQFJjsmcbipJgC2MpgQNTeczNg25CSeIWnboQqj6exQ
51fe6o/QPx8BL48BtM6+IS7yOkbGvdmf0ljDIzDX4KtoyL4c3cPhbwSEikxOMWwO
S1ta4eBD0HvjY2Scnmt2q887m2q0ICw0+wVn1XODrADP8Af+HSg/fJdPzDe3euaa
j8uXx4XNGBUloyiO9Tr1aIPB++1xYksgbUBwKRUi5rs7Hu9e0NnqlhLtc15tImUu
GnXu+9eFu+s+m06L2cZbFb2hYDrpzmHmLjLco5fW0503LzJwpIabNmtPcajJwgLX
8+74Ph+slnneXFmrYtgEmdB2fNEQ63pRjPPTYWAk+BSiHX58rJzcbLcQr6rLwnRM
4lG0sWZSVvpA1ndw5sWGmDU1aCt1j0EYwQZBRovJCThj6EI0+byJ9MnhtqgDx7nW
OElf4wGUPg1eF52W0S5HkDA53J6pzMfiFH6tXuKljWn6UmrofbyQKxrHj8RNtYJj
n0fi+1VOmW91T1hUcOF3Y9th1lvVApNi1hKNkwjsPDF7NV35CgjCGp0x9EoZS97w
jV4kOsl4cg1oJTyshTJNPr9m59E8UyydepSOjPNcvYIttOcpM4Z2uL1yy7LyF7AQ
uckWqTKUhkV2GhEFapAWYxwRspV4zCOehP07IUNGb73Z7AMnK9jN8O4m32RpLfIN
SQNaLFDu3WLWT6D28A1TUedkQXDawVHjYu4rDrKdul2iiDWpD/N0ODzL1ZRpMn5i
URqVm0rjUvowmw3bWMKQL9FN0znjvZ/TLLn/waqptQvAdsd6HNShc6giFEf0L7+4
UxC8seafJx4LZyEB5cBZd2vus56lftSLJ5qxoeFdfdjpzOk5ocJ3zDHGmg6zbENe
aYYoq6vZXBtlCOIIyI+Gkki4bSCmrYAC1CBIbEts5BWhQlytfuW5x7TF2mw0J4ZV
fYfUvBoIpMgyX7AQzNnzCeaDvKg82GICEoeCc6k037B/1VenJN1KocvD72Yn8QIY
ZS98ltabksOA7oWcY4RIhXqnmvNQVmhoPZTnkLR04Ey5PK8cqwteatZIIxp1T2gW
cGIdq1ToB92Pv17fhaKk8jaeWcWjLqV/co/W+LXBzZCKa9zM2EPOw9I3UDLzeixU
vuByI2wy7/YVnfEhRy1JNPFFqB23Yg+pZ4D7zWSeUDu9oT6q9MLeGuZO/aDkaIjh
v5R+uAgjwULQ9o5GJndaTNMfZ6yTgIqp2YT0JRUPq4Z9GGyatq+aMc9ADMFPYV7h
5wnhvKygHxeOBF13FSB4clG0mMH7II6EqABL+s5ugIjlYAJjpD+044a7BjpIr2A+
VcZo5hhK429poj3GFufbJX2WEEgQulqL1QqKwZw/OmoMTkHlzGRl/1dguqHKyE4r
5inxvJuqYym2prQgHr4HN/ucMhUqYdL1iN2zoE6Jh87GrQYS7kT9fs9x7orOchBI
iQE36OPFMTSsP+1CsGY3tnWA7zGOzhk1F1wCdfk1tIe60cUMLdcpZV0a6eWybV2w
zcvsddMNI2N2IvzSZ5WNysaldGDm+qNgU7pxrIhOZmSI1RQDzQSF8oFL5k2bQwtN
MuFojGJyRrPz01wm17U96IR0zpWlUnEXwZhDwoek9K4Kx3Q32tpsVpL2SUkIGKl7
pxWGjaW3DN4jzkiEB6DztpICiFV2Nkz3ThuKgNqgXJeLdgax0JBB6suBqbjjdCqh
sOkZKddL+ShfkiuN4wmzV1GJZpotNM5nAklItjQiI9SluHw4dZfhDz7APgKnRIw0
w9pdifDo/7/NLmqlinlEbBHZKz0KktTLBii8lkAUmaVhqZ6kp3UK1gQvMT8SsdSa
gYIMGsvoX6/4BzDEKKyaoay0DbJ9iAt0jRGNnbIr3ckSkxbmWkjcGemVmkHnY6FE
XxcoFh0CUQsYlQ+1hO8HmCHXt1TmAD03FgrOtP0jTm0UCXgv5Fh5FSmt06ZHa3WY
yiuD/r8LPSodlerYizPC/v0K0aiBGUbFkdvtoj4BP/DTM9V6QfUBYbchQ8LnoAzu
9YoCFiGlZfui5WyPjmT+OiQK+C23r3dHnAmayb9CA3RlEujfW1tWvrsUs17g97pH
Kw1p7g0x4CHFrgeytqZvTNQCA3Zxpy5y5cJ3LsEU+7F9yMfXiTESmVmz9wGbE2bp
d12/K3kLl0wx8ivF/bq/g5Z1JOHOL0O9ZcyqiXtH60HeCWzNaT6BB8gRZ7+QaULK
teRtqCH9zJDHFN4PH09LI+A2woJ+xCxLBM2KWzzez88g1UVDRXi4bAQp10Wz/dA9
0G5ypqebAXVv1H4luHPGPEiw6tx+ALXlTTgOPt/eDVQMbT2w6UdxUHwqEj+FNWgf
+xtwDfsQsJbnBqFXHicM46sepKCYP9iPCj6EOJrC1m9C8u0/Tp/QI2d1OcbjPldz
MxO+G5GVEF/w1A3adPwZJmdITxhhUtJl05fikAszyxE61sXTqu16FsZuuPx0o1Po
Kh35q3thvH2p5kCjoNUJsOekxLXEdsJeRz6C4oT9uzdCXWxktg7oHmtwy0qYdUV6
8azrtbto1RucCN+NuCR+QbVhwQLU52vHWRwR1ANE90NJ4OQdSToLMslU0FqNm5bP
8ND9/kMa6Q2qqgR8hvRHXye1M2ZOJ/+rRh0l1dw2J/pub5lYDLB+SfhSF90d0vck
Ku44XEVYij6o/57xm400aSWi0OnUYPLuhuIxidLzv54UMkN5BqOY2Cyby2G2CjJP
eDg3ATjHgg9ApTBS0/tlkRrD9VlH2gCwqV3LYroIDNgRwmZs/nwlZUQG4nzw6wYV
tTehvSAhA/+8bRtJQiobmveUA00XTpGQmU64rUxpLvHLlPrEvNN4k8ovTiuDte6a
y1iom323lqGtUo27ki4HbbiDVvZLHqHXQ4Q4roIDSzqc2Zw9E30cghc/s1T5thaH
TFiR7JKX1bzelG+yrCveMaCoui/yZRMLCJ5dXQDEytVuXTBJ9Pjr46iTnCOO22O/
ay/jgeddC+7hC3uH+8oMMvFXHraxSXM5zQgKuQ6Wgco89LZIf8v+BSDBsoFGlm3g
Q9FAKmUF5NgL91jqSVJt4fAfULrCAapKeGV/Z5KVxQ4tQ9CSbidec4AOwwG9s1up
80TCB8qpOSfAYhomGfHsLHgSLYQqx0xoU0I79hAGdshzg9zcjXKejJ6hSHGOW/Ph
0nK4TcR7tbxNt1/czvrJtjHC2h7qyglIe95H/voW34/S/wigyYa3SUb/c4Chxln9
v7cDBJEP6qZqbZI0rreZxl63NqPwH1Z40lAGehLBUrHQseEbyS/W3MX4jv6OCiys
KG/HX/Z6y6F1De052MnqjBzrYoKHySvxp67cTkhLGqeQr4yV2d4KX2162HF5rr4f
BCnliKpZKeWOG3SUNA1qpias5ViIDkaHopyfrpMF1/P7Rpt6O6391yQSDH2E6uj4
68St18APHR3W+T5nAUTAOocRlR9exWCvYUtt2i+TxnESe7yl8/bEY0KcQpdhxZ4Y
PB6Nm9X4StDoh34bOJ0Ye9rqwwLwBMntkIZJN12H9yN7iRNRqd79aQf9/SOZIyT/
5VsBY1V1xzgIjBMEZjYR4gs09AqpAy37dEoqLMFqCOTahFFH9jUmkLA0mCbRTKzR
G6ushfI/LpHZtnV9lVeSDzZTOfAZhKwFfwpwIh7SOcuzbmJtz6G0Ij7FCwRzfJjK
6wk5BVr88YcjnEVNSImz18wuwtkRH6CL/bcVzXGlJo+ThJ58Nqp6ElG7sMSwHav9
KIKqaszTKfiGSBRjbeF7yySIYB2T+wA3/Cs1S7EpDvhRLZSfaCRlWgoTdmLNCLeV
CBCvFox9rndyHOBjvHQD/HpWWi8Wm/l8OGQqyXkSka93VTGXxURnVRkqQWNnGsxk
yKcdhdyzE5yhFbwVVBecMhKGoqjrxUmNGe3ycJ/P/E6GA13vn9wSAXJHqf70K/07
A6qcUMWijdFdw7J0aD88YnQw7Jde42bA9YbnMdPF+8lQF27RS8DXRhkXL3NKoIHg
0ezauvJFb7gk5D5pVzWMkwgX8BMP+rNSmV5S/akxM6jY+LD4NB+SCwezMkLsBzQX
2ewOhGS8H8KnW3LIUvb784ssXo+9Vi04GRPmy0F4vzSSV8oLXArqELM5gw7RZjJE
x6Xsmi3I5nBEuEAZMlwS5+9sRhvWG8UrwnhhbokpE6ltaWDYKIzUFhKcXprgglpC
7xKCMEgo+Xx+NB2wkxFgmMiPIY5+N12dH4K6sroHiHwhzrMqOsen93CPsRZDs1m4
V5u4zWxYzhn1MVQDu9IuNvXir6juMaYxAd1ywfRQ6CyVcr5im0fGAxc7LmrGyJVO
zvgF7uzv27i4vRFU7G7UCaK1xmupXQTB29/pcDfpHTu8OWRc8+KQ1f8BEj/Tebi1
oELMV+YiGB7MgWLzPrGoVQNeSkhGO43GO2ou1ITtf3a1i5LY6CXwqpKmDnGvZD2z
fo6K7cuL302wnumdsHeto66S+rFmDs6krbmHshbaL5tnL94Q/x2q0Z+1nw1KfNJn
SNWapZ0nH/m65r6Nn/7cMVzgvPARwdjmKWWEuR96jekTY/UKTQJ/XqxDiaHSacjy
euFmzBDy3bvau8qBmPNO0irJhXV7PbUDlTCFM9qEEJXvpBm/wwDOK8WYOCrZNLrj
oOJJFE35EBrfGlUVT1PiF0gg9EU9+Vki70N43jIqQ0ErhtnzEzl3GaupBWPWFAr/
r1UVxnNBUX/f/SvOCZFg6tYt3FMaTf35CzvmjHsXqN/ioHTa3xBuYpAuUF1WP9V/
j78bY/s7gSjhezA4qnE+r0NEZBVfUu1i91/IyjGTH1is/Ka6NEPmR957ZmcVcQsn
QUpZ/PdD5yOko8BHPKl35Es59OPrxSfx2jNGeBkkGF4gidw5Fcq0MJB5TUAtjFQu
73Af1wmX3cRWLqTdSX1dyh0c2+gbzuXnqZ014AE08ojrWW3a29XLB/q9T2BsaM2r
7XUjeQPYutR60ZCycEmZZC11V/Jv4W05EFWx+U4WJ87+SGrlAGeu3qPJPFzh+pFe
Y8xbTCyV5CeJFJbayaXKah2Uh9LZTbf2BFpTqcGQv6ySGXMCWvO+sH7NwOkDF/gw
kEe45EsEiQfUWKkBggLCzO3PZkafcbPQl6/Agt6GArXqWiyD+krO5YD/3m93v4vY
ZLCl6807mzBIAvnBWt63fDzL3jt6JLkvRbQVjao2cr1f3gfzvhTegVX18k8eTnKa
j3ioj2gJEMIk/+Z9X/9tkzinhWjMxx1XGSeWhIp7KZFnBB4tWDm3F0Zx09bBsGgF
L/95Od7PPzX8Sy55auL8OcpFevh8dtzD/mjVgTdC/i79GVLDkV7hp/X+PP17OWLk
PcI8YNwdNwq1X790tDIdpG5kizwISSc/qbJKZhRRfjtwD5IC1a8txwpXdJTeoRLk
NikSRVZ9WdyfWVRteWyfUaJjCDOCH/nvGhZBuhrV84VmA5AVQIJeBkyMmeA72EV1
H0Z8bl+eXtmyfXSvtVSP7fHvrly2QVpQwO++EKJhCoXSIca8/z3yYc0l74pfpLLB
nZTB5PgGpsetiP2ZaBM0vYKxrpvTjTPDL0Vp2vJrJ8wgjWoiKqdMjRFGe0042P4d
OW0wyvWJN8tJ8HXaKu5NZlNnlvVjyyXSY43m6YxFrBffd63X21kOLCcvi2/EfQDa
zbj9va4a7MCW0WTNWWVav6pzXJTHOrEuSeYQ9HhJwPqWraUYfdgcowNJbior4fv9
oN6SXM9fGY6r5PX2/8Irt1tMtvYdO6HkqLkXHMyScrcHgPfmm1YBljttpCUwqiLS
k6zMn7o8vppUE9b9LWJErF1vHeVTEZU0vcjpdWrGyrWuGXlngnJP1ta7ssSj99uc
NqhegTABhhd8L1nVuy203hrmQSomn1ohfo6yhHUCcRbCZWuAUL9mNafIRzGxMNG5
5TpKPyC8VZJSMu/1k2nJ3S4g9DCqwgGQcnRwuvrIEob+HRkhuQSwZ3mdv5VN1sQV
JuWW8nrZU3TjgSyNtxZqetpN/6aNBsEdSKhaED1oiXWL8DpV5cbRvLyvOMBn+e3r
P8rF9hzZXU5D3cxWUocJ0s29++6PsPLIsyLhngKpXOKEmzIdNjIk29XNYYeOmPXI
J+yjgqp/b1iyvlzBDJlDMAM+uhjRs6b+Jl3PAHbC7NjxPQjJdcFL1wrBLF2jOXF6
F1y9QTPhc0+CVqyqSsZpD+aETd7ijXcHIuPGj0VALg649ixgrw98XCOsNAKwgTJh
5CthtQYENJ6r8k2VCenuRlIjm9LzE/NwiGhTaPZmApxuS2r7CH9cTa1LjoxFl/7w
8pIkywQQiKGvlJW0wHE0sURlRFmzVqsLl9HtHrHqnB616eBSxO3xMl0bFi5znlre
NNxHUsUBsyDdAA1EjMKgq3UpCe+tCLwLL8UpC7NRyMaKyKNtSTQ+JpUlp6Y0g8AZ
zWUlUuIiAFoSWX5fqocSUllnCvRRsLwTIKgueCJM6kYtUsr6FV1vrpP31Kk4Sywc
KguWq7xiPlHHTgcetCJL2co/kb6c68DFkZNhBlqs7itaI4irXzE44kYgi1hfYKxy
xxhpeu2HUVotrox5q3JOA11xm79wJDZZIg/izUP002XwVT/7U3HWN0/Wu+jl/Aa6
Rg1TNlwX8Mbqv4DWYLV+jxlo6sLrLSP7+b14Vh0Hf8JtLJjA7kAD+WUPpDA+V1kS
cSNWS72jZqJimep5YHjETbjEt/XSa7ENqBsV1bSegXg8aLaqoRhNe6YpQFVK2M/J
SEZpUErwgTBg4/g2kxodieu69TYSxv4UQUSaprY+I+xnaESb/1gehCasuKrdKuj9
D79DghjzroCFrZFaYfwAWHt7VYbAsB0rscsLzFpxagUEXwk/6tb9X2pOk70jNja7
//H6zr51qOda6rNPuaMBiBkEvmaFkN3CVZy3g0r1macZPjqa72rnSd94+EjSHpum
upushTXTGnaK71WFEA/2X0WYYN+7/DQ8EOnaFSY/ATgBNlLK0aFYXfXC4cSSTE+9
J5ShjlFTfsbPP1bD73uj6SJTMHdDnJG0nnlQl/5EjD8JZ33ab3XB2Mn5SxE1g6oq
uNTPpC2bVWzQgayivX02oZGSQ56HBBinXZXPcHbaJGn5CgWM/UrX2aQ68nERhCzz
EBGwIwUvcIIuIYR2AQso2ctyzYQQyZRRlZOnmEqvNKkf9KTHlYB5teHwA1DC9/zf
duYKh//bRIqRwdJip0uaJ3FapjDVrpboPNRWBjwjCpimdDNFnUnwAfPYbKSKS1fu
K35DTR+dQt4BxDVTF+yVZcL7LP+MeYGRERvJcnkUVrLAWg6eywyPN/C9BvW8COzV
ghcsFgN2kNE9iO2dTQPE7arIVVI31cGSxA3AFQ6mdOWlkuc9RgfnQm0AltAnSQqV
pWhLXxlCnZCYR4koP9+7opp2Y9qUlw8/wUef/zG1CsoRouBRUlnmf39AUSAa+xbT
H//0c56GZBdbjT25q3XmpA6xDQ+RK8F+VikwBtIbc7R3U+0U2RhAjx58h2yVtlPO
CYdnwU7KqhPNCExRtuRasX0Eg4vdGSGz26d7wsDk5yu576KTLWW4VMs6awqXGa10
C2pWmYfkfVg360ZkpVnzGp9Q3eDVCKQ4ardS0r5TsKu8Mu+z4QVUwxUCe6uzgBZr
4MxXt2Bye98t1L1Ig18fFJ7AAmpNVt8X1PXmWEVqbz3QugBa5srCousArYLlyTB4
+gdKrw4UdeTzYhtsjuHXqbw/xuUg5nUNk2tvrQV2JsBPoiOz0BW1yH1HUSv7lcCd
jGn34Gkz5ld+Rqyct0wmeZhzBNXxKbqZ1IgKIQXtlX4n7hRL6dr6LRQz4ToxZw2N
FGIvCn2vU87u9Hg95e4Psu++uYZ/uoKGCSNO021bh9VEaVvEZQGZ94HEugT/hk1t
r9Sw2ac8Sd9qRyN7wasGEPoU3Pd7zgGWvkimrS/zWEPbb7F5kixA3SXTfHM4sWPH
1h2dObznAuqvLcMKWeONV2XISNR1rDuGJ2a8iN+AHN9DAW+ZBpkNyKG3X+2aer0V
xCPPgbNBUp3oXG7sJmc7NooIkKfMBPfMgsk7RzsgQRY386TD+BSCeoJFsl9jl7Yt
Ic+FN71rTeHVgJ8+UM10m1ldKGqiX57sIDK7KbsvraJU1wUBYS5UnbRHXeNBVGRW
1BiFvtJNi/mnxi+QYCr78qAQNIVopb2LkYhS4iLIeFxYJfEln6PgwuWnJRrq+Icj
4IqsluGlPrBDjuwfbxWBm2DgFtsb3XO4tESu+mGG1AIMux1mfrcVqzNnqj+izysg
kVTyIH228Wt/MH8a4/VRsw==
//pragma protect end_data_block
//pragma protect digest_block
W7qLMrdCsI4q9lhFda8Pqh78/0M=
//pragma protect end_digest_block
//pragma protect end_protected
